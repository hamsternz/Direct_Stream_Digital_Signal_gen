library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

entity dsdsg is
   port ( clk100MHz : in  std_logic;
          pin       : out std_logic);
end entity;

architecture whatever of dsdsg is
  signal addr : unsigned(11 downto 0) := (others => '0');
  signal data : std_logic_vector(31 downto 0) := ( 0 => '1', others => '0');
  signal mask : std_logic_vector(31 downto 0) := ( 0 => '1', others => '0');
  type a_memory is array (0 to 3124) of std_logic_vector(31 downto 0);
  signal memory : a_memory := (
     "10101010101010101010101010101010",  --  0.0000000 -  0.0019478
     "10101010101010101010101010101010",  --  0.0020106 -  0.0039584
     "10101010101010101010101010101010",  --  0.0040212 -  0.0059690
     "10101010101010101010101010101010",  --  0.0060319 -  0.0079796
     "10101010101010101010101010101010",  --  0.0080425 -  0.0099903
     "10101010101010101010101010101010",  --  0.0100531 -  0.0120009
     "10101010101010101010101010110101",  --  0.0120637 -  0.0140115
     "01010101010101010101010101010101",  --  0.0140743 -  0.0160221
     "01010101010101010101010101010101",  --  0.0160850 -  0.0180327
     "01010101010101010101011010101010",  --  0.0180956 -  0.0200434
     "10101010101010101010101010101010",  --  0.0201062 -  0.0220540
     "10101010101010101010101010110101",  --  0.0221168 -  0.0240646
     "01010101010101010101010101010101",  --  0.0241274 -  0.0260752
     "01010101010101010101011010101010",  --  0.0261381 -  0.0280858
     "10101010101010101010101010101010",  --  0.0281487 -  0.0300965
     "10101010101101010101010101010101",  --  0.0301593 -  0.0321071
     "01010101010101010101010110101010",  --  0.0321699 -  0.0341177
     "10101010101010101010101010101010",  --  0.0341805 -  0.0361283
     "10101101010101010101010101010101",  --  0.0361911 -  0.0381389
     "01010101010110101010101010101010",  --  0.0382018 -  0.0401496
     "10101010101010101101010101010101",  --  0.0402124 -  0.0421602
     "01010101010101010101011010101010",  --  0.0422230 -  0.0441708
     "10101010101010101010101101010101",  --  0.0442336 -  0.0461814
     "01010101010101010101010110101010",  --  0.0462442 -  0.0481920
     "10101010101010101010101101010101",  --  0.0482549 -  0.0502027
     "01010101010101010101101010101010",  --  0.0502655 -  0.0522133
     "10101010101010101101010101010101",  --  0.0522761 -  0.0542239
     "01010101010110101010101010101010",  --  0.0542867 -  0.0562345
     "10101011010101010101010101010101",  --  0.0562973 -  0.0582451
     "01101010101010101010101010110101",  --  0.0583080 -  0.0602557
     "01010101010101010101101010101010",  --  0.0603186 -  0.0622664
     "10101010101011010101010101010101",  --  0.0623292 -  0.0642770
     "01011010101010101010101010110101",  --  0.0643398 -  0.0662876
     "01010101010101010110101010101010",  --  0.0663504 -  0.0682982
     "10101011010101010101010101010110",  --  0.0683611 -  0.0703088
     "10101010101010101011010101010101",  --  0.0703717 -  0.0723195
     "01010101101010101010101010101101",  --  0.0723823 -  0.0743301
     "01010101010101011010101010101010",  --  0.0743929 -  0.0763407
     "10101101010101010101010110101010",  --  0.0764035 -  0.0783513
     "10101010101101010101010101010110",  --  0.0784142 -  0.0803619
     "10101010101010101101010101010101",  --  0.0804248 -  0.0823726
     "01011010101010101010110101010101",  --  0.0824354 -  0.0843832
     "01010110101010101010101011010101",  --  0.0844460 -  0.0863938
     "01010101011010101010101010110101",  --  0.0864566 -  0.0884044
     "01010101010110101010101010101101",  --  0.0884672 -  0.0904150
     "01010101010101101010101010101011",  --  0.0904779 -  0.0924257
     "01010101010101101010101010101011",  --  0.0924885 -  0.0944363
     "01010101010101101010101010101011",  --  0.0944991 -  0.0964469
     "01010101010101101010101010101101",  --  0.0965097 -  0.0984575
     "01010101010110101010101010110101",  --  0.0985203 -  0.1004681
     "01010101011010101010101011010101",  --  0.1005310 -  0.1024788
     "01010101101010101010101101010101",  --  0.1025416 -  0.1044894
     "01010110101010101011010101010101",  --  0.1045522 -  0.1065000
     "01101010101010110101010101010110",  --  0.1065628 -  0.1085106
     "10101010101101010101010101101010",  --  0.1085734 -  0.1105212
     "10101011010101010101101010101010",  --  0.1105841 -  0.1125318
     "10110101010101011010101010101101",  --  0.1125947 -  0.1145425
     "01010101011010101010101101010101",  --  0.1146053 -  0.1165531
     "01011010101010101101010101010110",  --  0.1166159 -  0.1185637
     "10101010101101010101011010101010",  --  0.1186265 -  0.1205743
     "10110101010101011010101010101101",  --  0.1206372 -  0.1225849
     "01010101101010101010110101010101",  --  0.1226478 -  0.1245956
     "10101010101011010101010110101010",  --  0.1246584 -  0.1266062
     "10101101010101011010101010101101",  --  0.1266690 -  0.1286168
     "01010101101010101011010101010101",  --  0.1286796 -  0.1306274
     "10101010101101010101011010101010",  --  0.1306903 -  0.1326380
     "11010101010101101010101011010101",  --  0.1327009 -  0.1346487
     "01011010101010110101010101101010",  --  0.1347115 -  0.1366593
     "10101101010101011010101010110101",  --  0.1367221 -  0.1386699
     "01010110101010101101010101011010",  --  0.1387327 -  0.1406805
     "10101011010101011010101010110101",  --  0.1407434 -  0.1426911
     "01010110101010101101010101011010",  --  0.1427540 -  0.1447018
     "10101101010101011010101010110101",  --  0.1447646 -  0.1467124
     "01011010101010110101010101101010",  --  0.1467752 -  0.1487230
     "10110101010101101010101101010101",  --  0.1487858 -  0.1507336
     "01101010101101010101011010101011",  --  0.1507964 -  0.1527442
     "01010101011010101011010101010110",  --  0.1528071 -  0.1547549
     "10101011010101011010101010110101",  --  0.1548177 -  0.1567655
     "01011010101011010101010110101010",  --  0.1568283 -  0.1587761
     "11010101011010101011010101010110",  --  0.1588389 -  0.1607867
     "10101011010101011010101011010101",  --  0.1608495 -  0.1627973
     "01101010101101010101101010101011",  --  0.1628602 -  0.1648080
     "01010101101010101101010101101010",  --  0.1648708 -  0.1668186
     "10110101010110101010110101010110",  --  0.1668814 -  0.1688292
     "10101011010101011010101011010101",  --  0.1688920 -  0.1708398
     "01101010101101010110101010110101",  --  0.1709026 -  0.1728504
     "01011010101011010101011010101011",  --  0.1729133 -  0.1748610
     "01010101101010110101010110101010",  --  0.1749239 -  0.1768717
     "11010101011010101011010101101010",  --  0.1769345 -  0.1788823
     "10110101010110101011010101011010",  --  0.1789451 -  0.1808929
     "10101101010101101010110101010110",  --  0.1809557 -  0.1829035
     "10101101010101101010101101010110",  --  0.1829664 -  0.1849141
     "10101011010101101010101101010101",  --  0.1849770 -  0.1869248
     "10101011010101011010101101010101",  --  0.1869876 -  0.1889354
     "10101011010101011010101101010101",  --  0.1889982 -  0.1909460
     "10101011010101011010101101010101",  --  0.1910088 -  0.1929566
     "10101011010101101010101101010110",  --  0.1930195 -  0.1949672
     "10101011010101101010110101010110",  --  0.1950301 -  0.1969779
     "10101101010110101010110101011010",  --  0.1970407 -  0.1989885
     "10110101010110101011010101101010",  --  0.1990513 -  0.2009991
     "11010101011010101101010110101011",  --  0.2010619 -  0.2030097
     "01010101101010110101011010101101",  --  0.2030725 -  0.2050203
     "01011010101011010101101010110101",  --  0.2050832 -  0.2070310
     "01101010110101011010101011010101",  --  0.2070938 -  0.2090416
     "10101011010101101010110101011010",  --  0.2091044 -  0.2110522
     "10110101011010101101010101101010",  --  0.2111150 -  0.2130628
     "11010101101010110101011010101101",  --  0.2131256 -  0.2150734
     "01011010101101010110101011010101",  --  0.2151363 -  0.2170841
     "10101011010101101010110101011010",  --  0.2171469 -  0.2190947
     "10110101011010101101010110101011",  --  0.2191575 -  0.2211053
     "01011010101101010110101011010101",  --  0.2211681 -  0.2231159
     "10101011010101101010110101011010",  --  0.2231787 -  0.2251265
     "10110101101010110101011010101101",  --  0.2251894 -  0.2271371
     "01011010101101010110101101010110",  --  0.2272000 -  0.2291478
     "10101101010110101011010110101011",  --  0.2292106 -  0.2311584
     "01010110101011010101101011010101",  --  0.2312212 -  0.2331690
     "10101011010101101011010101101010",  --  0.2332318 -  0.2351796
     "11010101101011010101101010110101",  --  0.2352425 -  0.2371902
     "10101011010101101011010101101010",  --  0.2372531 -  0.2392009
     "11010110101011010101101011010101",  --  0.2392637 -  0.2412115
     "10101011010110101011010101101011",  --  0.2412743 -  0.2432221
     "01010110101011010110101011010110",  --  0.2432849 -  0.2452327
     "10101101010110101101010110101101",  --  0.2452956 -  0.2472433
     "01011010101101011010101101011010",  --  0.2473062 -  0.2492540
     "10110101101010110101101010110101",  --  0.2493168 -  0.2512646
     "10101011010110101011010101101011",  --  0.2513274 -  0.2532752
     "01010110101101010110101101010110",  --  0.2533380 -  0.2552858
     "10110101101010110101101010110101",  --  0.2553487 -  0.2572964
     "10101011010110101011010110101011",  --  0.2573593 -  0.2593071
     "01011010110101011010110101011010",  --  0.2593699 -  0.2613177
     "11010101101011010110101011010110",  --  0.2613805 -  0.2633283
     "10101101011010110101011010110101",  --  0.2633911 -  0.2653389
     "10101011010110101011010110101101",  --  0.2654017 -  0.2673495
     "01011010110101101010110101101011",  --  0.2674124 -  0.2693602
     "01010110101101011010101101011010",  --  0.2694230 -  0.2713708
     "11010101101011010110101101010110",  --  0.2714336 -  0.2733814
     "10110101101010110101101011010110",  --  0.2734442 -  0.2753920
     "10101101011010110101101010110101",  --  0.2754548 -  0.2774026
     "10101101011010101101011010110101",  --  0.2774655 -  0.2794133
     "10101011010110101101011010101101",  --  0.2794761 -  0.2814239
     "01101011010110101101010110101101",  --  0.2814867 -  0.2834345
     "01101011010110101101010110101101",  --  0.2834973 -  0.2854451
     "01101011010110101011010110101101",  --  0.2855079 -  0.2874557
     "01101011010110101101010110101101",  --  0.2875186 -  0.2894663
     "01101011010110101101011010101101",  --  0.2895292 -  0.2914770
     "01101011010110101101011010110101",  --  0.2915398 -  0.2934876
     "10101101010110101101011010110101",  --  0.2935504 -  0.2954982
     "10101101011010110101101011010110",  --  0.2955610 -  0.2975088
     "10110101101010110101101011010110",  --  0.2975717 -  0.2995194
     "10110101101011010110101101011010",  --  0.2995823 -  0.3015301
     "11010110101101011010110101101011",  --  0.3015929 -  0.3035407
     "01011010110101101011010110101101",  --  0.3036035 -  0.3055513
     "01101011010110101101011010110101",  --  0.3056141 -  0.3075619
     "10101101011010110101101011010110",  --  0.3076248 -  0.3095725
     "10110101101011010110101101011010",  --  0.3096354 -  0.3115832
     "11010110101101011010110101101011",  --  0.3116460 -  0.3135938
     "01101011010110101101011010110101",  --  0.3136566 -  0.3156044
     "10101101011010110101101011010110",  --  0.3156672 -  0.3176150
     "10110110101101011010110101101011",  --  0.3176778 -  0.3196256
     "01011010110101101101011010110101",  --  0.3196885 -  0.3216363
     "10101101011010110101101011011010",  --  0.3216991 -  0.3236469
     "11010110101101011010110101101101",  --  0.3237097 -  0.3256575
     "01101011010110101101011010110110",  --  0.3257203 -  0.3276681
     "10110101101011010110101101101011",  --  0.3277309 -  0.3296787
     "01011010110101101101011010110101",  --  0.3297416 -  0.3316894
     "10101101011011010110101101011010",  --  0.3317522 -  0.3337000
     "11011010110101101011010110110101",  --  0.3337628 -  0.3357106
     "10101101011011010110101101011010",  --  0.3357734 -  0.3377212
     "11011010110101101011011010110101",  --  0.3377840 -  0.3397318
     "10101101101011010110101101101011",  --  0.3397947 -  0.3417424
     "01011010110110101101011010110110",  --  0.3418053 -  0.3437531
     "10110101101011011010110101101011",  --  0.3438159 -  0.3457637
     "01101011010110110101101011010110",  --  0.3458265 -  0.3477743
     "11010110101101101011010110110101",  --  0.3478371 -  0.3497849
     "10101101011011010110101101101011",  --  0.3498478 -  0.3517955
     "01011011010110101101101011010110",  --  0.3518584 -  0.3538062
     "11010110101101101011010110110101",  --  0.3538690 -  0.3558168
     "10101101101011010110110101101011",  --  0.3558796 -  0.3578274
     "01101011010110110101101011011010",  --  0.3578902 -  0.3598380
     "11011010110101101101011010110110",  --  0.3599009 -  0.3618486
     "10110101101101011011010110101101",  --  0.3619115 -  0.3638593
     "10101101101011010110110101101011",  --  0.3639221 -  0.3658699
     "01101011011010110101101101011011",  --  0.3659327 -  0.3678805
     "01011010110110101101101011011010",  --  0.3679433 -  0.3698911
     "11010110110101101101011011010110",  --  0.3699540 -  0.3719017
     "10110110101101101011011010110101",  --  0.3719646 -  0.3739124
     "10110101101101011011010110101101",  --  0.3739752 -  0.3759230
     "10101101101011011010110110101101",  --  0.3759858 -  0.3779336
     "10101101011011010110110101101101",  --  0.3779964 -  0.3799442
     "01101101011011010110110101101101",  --  0.3800070 -  0.3819548
     "01101101011011010110110101101011",  --  0.3820177 -  0.3839655
     "01101011011010110110101101101011",  --  0.3840283 -  0.3859761
     "01101011011010110110101101101011",  --  0.3860389 -  0.3879867
     "01101011011011010110110101101101",  --  0.3880495 -  0.3899973
     "01101101011011010110110101101101",  --  0.3900601 -  0.3920079
     "01101101011011010110110110101101",  --  0.3920708 -  0.3940186
     "10101101101011011010110110101101",  --  0.3940814 -  0.3960292
     "10101101101101011011010110110101",  --  0.3960920 -  0.3980398
     "10110101101101101011011010110110",  --  0.3981026 -  0.4000504
     "10110110110101101101011011010110",  --  0.4001132 -  0.4020610
     "11011010110110101101101011011011",  --  0.4021239 -  0.4040716
     "01011011010110110110101101101011",  --  0.4041345 -  0.4060823
     "01101101011011010110110110101101",  --  0.4061451 -  0.4080929
     "10101101101101011011010110110110",  --  0.4081557 -  0.4101035
     "10110110101101101101011011010110",  --  0.4101663 -  0.4121141
     "11011010110110110101101101011011",  --  0.4121770 -  0.4141247
     "01101011011011010110110110101101",  --  0.4141876 -  0.4161354
     "10101101101101011011011010110110",  --  0.4161982 -  0.4181460
     "11010110110110101101101011011011",  --  0.4182088 -  0.4201566
     "01011011011010110110110101101101",  --  0.4202194 -  0.4221672
     "10101101101101011011011010110110",  --  0.4222301 -  0.4241778
     "11010110110110101101101101011011",  --  0.4242407 -  0.4261885
     "01101011011011010110110110110101",  --  0.4262513 -  0.4281991
     "10110110101101101101011011011010",  --  0.4282619 -  0.4302097
     "11011011011010110110110101101101",  --  0.4302725 -  0.4322203
     "10101101101101101011011011010110",  --  0.4322831 -  0.4342309
     "11011011010110110110101101101101",  --  0.4342938 -  0.4362416
     "10101101101101011011011011010110",  --  0.4363044 -  0.4382522
     "11011010110110110110101101101101",  --  0.4383150 -  0.4402628
     "10101101101101101011011011010110",  --  0.4403256 -  0.4422734
     "11011011010110110110110101101101",  --  0.4423362 -  0.4442840
     "10110101101101101101011011011011",  --  0.4443469 -  0.4462947
     "01011011011011010110110110110110",  --  0.4463575 -  0.4483053
     "10110110110110101101101101101011",  --  0.4483681 -  0.4503159
     "01101101101011011011011011010110",  --  0.4503787 -  0.4523265
     "11011011010110110110110110101101",  --  0.4523893 -  0.4543371
     "10110110110101101101101101011011",  --  0.4544000 -  0.4563477
     "01101101101011011011011011010110",  --  0.4564106 -  0.4583584
     "11011011011010110110110110110101",  --  0.4584212 -  0.4603690
     "10110110110110101101101101101101",  --  0.4604318 -  0.4623796
     "01101101101101101101011011011011",  --  0.4624424 -  0.4643902
     "01101011011011011011011010110110",  --  0.4644531 -  0.4664008
     "11011011011010110110110110110110",  --  0.4664637 -  0.4684115
     "10110110110110110110101101101101",  --  0.4684743 -  0.4704221
     "10110110101101101101101101101011",  --  0.4704849 -  0.4724327
     "01101101101101101101011011011011",  --  0.4724955 -  0.4744433
     "01101101011011011011011011011010",  --  0.4745062 -  0.4764539
     "11011011011011011011011010110110",  --  0.4765168 -  0.4784646
     "11011011011011010110110110110110",  --  0.4785274 -  0.4804752
     "11011011010110110110110110110110",  --  0.4805380 -  0.4824858
     "11010110110110110110110110110101",  --  0.4825486 -  0.4844964
     "10110110110110110110110110101101",  --  0.4845593 -  0.4865070
     "10110110110110110110110101101101",  --  0.4865699 -  0.4885177
     "10110110110110110110110101101101",  --  0.4885805 -  0.4905283
     "10110110110110110110110101101101",  --  0.4905911 -  0.4925389
     "10110110110110110110110110101101",  --  0.4926017 -  0.4945495
     "10110110110110110110110110110110",  --  0.4946123 -  0.4965601
     "10110110110110110110110110110110",  --  0.4966230 -  0.4985708
     "11011011010110110110110110110110",  --  0.4986336 -  0.5005814
     "11011011011011011011010110110110",  --  0.5006442 -  0.5025920
     "11011011011011011011011011011011",  --  0.5026548 -  0.5046026
     "01101101101011011011011011011011",  --  0.5046654 -  0.5066132
     "01101101101101101101101101101101",  --  0.5066761 -  0.5086239
     "10110110101101101101101101101101",  --  0.5086867 -  0.5106345
     "10110110110110110110110110110110",  --  0.5106973 -  0.5126451
     "11011011011011011011011010110110",  --  0.5127079 -  0.5146557
     "11011011011011011011011011011011",  --  0.5147185 -  0.5166663
     "01101101101101101101101101101101",  --  0.5167292 -  0.5186769
     "10110110110110110110110110110110",  --  0.5187398 -  0.5206876
     "11011011011011011011011011011011",  --  0.5207504 -  0.5226982
     "01101101101101101101101101101101",  --  0.5227610 -  0.5247088
     "10110110110110110110110110110110",  --  0.5247716 -  0.5267194
     "11011011011011011011011011011011",  --  0.5267823 -  0.5287300
     "01101101101101101101101101101101",  --  0.5287929 -  0.5307407
     "10110110110110110110110110110110",  --  0.5308035 -  0.5327513
     "11011011011011011011011011011011",  --  0.5328141 -  0.5347619
     "01101101101101101101101101101101",  --  0.5348247 -  0.5367725
     "10110110110110111011011011011011",  --  0.5368354 -  0.5387831
     "01101101101101101101101101101101",  --  0.5388460 -  0.5407938
     "10110110110110110110110110110110",  --  0.5408566 -  0.5428044
     "11101101101101101101101101101101",  --  0.5428672 -  0.5448150
     "10110110110110110110110110110111",  --  0.5448778 -  0.5468256
     "01101101101101101101101101101101",  --  0.5468884 -  0.5488362
     "10110110110110110111011011011011",  --  0.5488991 -  0.5508469
     "01101101101101101101101101101101",  --  0.5509097 -  0.5528575
     "11011011011011011011011011011011",  --  0.5529203 -  0.5548681
     "01101101110110110110110110110110",  --  0.5549309 -  0.5568787
     "11011011011011011101101101101101",  --  0.5569415 -  0.5588893
     "10110110110110110111011011011011",  --  0.5589522 -  0.5609000
     "01101101101101101101110110110110",  --  0.5609628 -  0.5629106
     "11011011011011011011101101101101",  --  0.5629734 -  0.5649212
     "10110110110110110111011011011011",  --  0.5649840 -  0.5669318
     "01101101101101110110110110110110",  --  0.5669946 -  0.5689424
     "11011011011101101101101101101101",  --  0.5690053 -  0.5709530
     "10111011011011011011011011011011",  --  0.5710159 -  0.5729637
     "10110110110110110110111011011011",  --  0.5730265 -  0.5749743
     "01101101101101110110110110110110",  --  0.5750371 -  0.5769849
     "11011101101101101101101101101110",  --  0.5770477 -  0.5789955
     "11011011011011011011101101101101",  --  0.5790584 -  0.5810061
     "10110110111011011011011011011101",  --  0.5810690 -  0.5830168
     "10110110110110110111011011011011",  --  0.5830796 -  0.5850274
     "01101110110110110110110111011011",  --  0.5850902 -  0.5870380
     "01101101101110110110110110110111",  --  0.5871008 -  0.5890486
     "01101101101101101110110110110110",  --  0.5891115 -  0.5910592
     "11011101101101101101101110110110",  --  0.5911221 -  0.5930699
     "11011011101101101101101101110110",  --  0.5931327 -  0.5950805
     "11011011011101101101101101110110",  --  0.5951433 -  0.5970911
     "11011011011101101101101101101110",  --  0.5971539 -  0.5991017
     "11011011011011101101101101101110",  --  0.5991646 -  0.6011123
     "11011011011011101101101101110110",  --  0.6011752 -  0.6031230
     "11011011011101101101101101110110",  --  0.6031858 -  0.6051336
     "11011011011101101101101110110110",  --  0.6051964 -  0.6071442
     "11011011101101101101110110110110",  --  0.6072070 -  0.6091548
     "11011101101101101110110110110111",  --  0.6092176 -  0.6111654
     "01101101101101110110110110111011",  --  0.6112283 -  0.6131761
     "01101101110110110110111011011011",  --  0.6132389 -  0.6151867
     "01101110110110110111011011011011",  --  0.6152495 -  0.6171973
     "10110110110111011011011011101101",  --  0.6172601 -  0.6192079
     "10110111011011011101101101101110",  --  0.6192707 -  0.6212185
     "11011011011101101101101110110110",  --  0.6212814 -  0.6232292
     "11011101101101101110110110111011",  --  0.6232920 -  0.6252398
     "01101101110110110110111011011011",  --  0.6253026 -  0.6272504
     "10110110110111011011011101101101",  --  0.6273132 -  0.6292610
     "10111011011011101101101101110110",  --  0.6293238 -  0.6312716
     "11011101101101101110110110111011",  --  0.6313345 -  0.6332822
     "01101101110110110111011011011101",  --  0.6333451 -  0.6352929
     "10110110111011011011101101101110",  --  0.6353557 -  0.6373035
     "11011011101101101101110110110111",  --  0.6373663 -  0.6393141
     "01101101110110110111011011011101",  --  0.6393769 -  0.6413247
     "10110110111011011011101101101110",  --  0.6413876 -  0.6433353
     "11011011101101101110110110111011",  --  0.6433982 -  0.6453460
     "01101110110110111011011011101101",  --  0.6454088 -  0.6473566
     "10111011011011101101101110110110",  --  0.6474194 -  0.6493672
     "11101101101110110110111011011011",  --  0.6494300 -  0.6513778
     "10110111011011011101101101110110",  --  0.6514407 -  0.6533884
     "11011101101101110110110111011011",  --  0.6534513 -  0.6553991
     "10110110111011011011101101101110",  --  0.6554619 -  0.6574097
     "11011101101101110110110111011011",  --  0.6574725 -  0.6594203
     "01110110111011011011101101101110",  --  0.6594831 -  0.6614309
     "11011101101101110110111011011011",  --  0.6614937 -  0.6634415
     "10110110111011011101101101110110",  --  0.6635044 -  0.6654522
     "11101101101110110111011011011101",  --  0.6655150 -  0.6674628
     "10110111011011101101101110110111",  --  0.6675256 -  0.6694734
     "01101101110110111011011011101101",  --  0.6695362 -  0.6714840
     "11011011101101101110110111011011",  --  0.6715468 -  0.6734946
     "01110110111011011101101101110110",  --  0.6735575 -  0.6755053
     "11101101101110110111011011101101",  --  0.6755681 -  0.6775159
     "10111011011101101110110110111011",  --  0.6775787 -  0.6795265
     "01110110111011011011101101110110",  --  0.6795893 -  0.6815371
     "11101101110110110111011011101101",  --  0.6815999 -  0.6835477
     "11011011011101101110110111011011",  --  0.6836106 -  0.6855583
     "10110111011011011101101110110111",  --  0.6856212 -  0.6875690
     "01101110110111011011011101101110",  --  0.6876318 -  0.6895796
     "11011101101110110111011011101101",  --  0.6896424 -  0.6915902
     "11011011011101101110110111011011",  --  0.6916530 -  0.6936008
     "10110111011011101101110110111011",  --  0.6936637 -  0.6956114
     "01110110111011011011101101110110",  --  0.6956743 -  0.6976221
     "11101101110110111011011101101110",  --  0.6976849 -  0.6996327
     "11011101101110110111011011101101",  --  0.6996955 -  0.7016433
     "11011011101101110110111011011101",  --  0.7017061 -  0.7036539
     "10111011011101101110110111011011",  --  0.7037168 -  0.7056645
     "10110111011011101110110111011011",  --  0.7057274 -  0.7076752
     "10110111011011101101110110111011",  --  0.7077380 -  0.7096858
     "01110110111011011101101110111011",  --  0.7097486 -  0.7116964
     "01110110111011011101101110110111",  --  0.7117592 -  0.7137070
     "01101110110111011101101110110111",  --  0.7137699 -  0.7157176
     "01101110110111011011101110110111",  --  0.7157805 -  0.7177283
     "01101110110111011011101110110111",  --  0.7177911 -  0.7197389
     "01101110110111011011101110110111",  --  0.7198017 -  0.7217495
     "01101110110111011101101110110111",  --  0.7218123 -  0.7237601
     "01101110110111011101101110110111",  --  0.7238229 -  0.7257707
     "01101110111011011101101110111011",  --  0.7258336 -  0.7277814
     "01110110111011011101110110111011",  --  0.7278442 -  0.7297920
     "01110111011011101101110111011011",  --  0.7298548 -  0.7318026
     "10110111011101101110110111011101",  --  0.7318654 -  0.7338132
     "10111011011101110110111011011101",  --  0.7338760 -  0.7358238
     "11011011101101110111011011101101",  --  0.7358867 -  0.7378345
     "11011101101110111011011101101110",  --  0.7378973 -  0.7398451
     "11101101110111011011101101110111",  --  0.7399079 -  0.7418557
     "01101110111011011101101110111011",  --  0.7419185 -  0.7438663
     "01110111011011101101110111011011",  --  0.7439291 -  0.7458769
     "10111011011101110110111011101101",  --  0.7459398 -  0.7478875
     "11011011101110110111011101101110",  --  0.7479504 -  0.7498982
     "11101101110111011011101110110111",  --  0.7499610 -  0.7519088
     "01110110111011101101110111011011",  --  0.7519716 -  0.7539194
     "10111011011101110110111011101101",  --  0.7539822 -  0.7559300
     "11011101101110111011011101110110",  --  0.7559929 -  0.7579406
     "11101110110111011101101110111011",  --  0.7580035 -  0.7599513
     "10110111011101101110111011011101",  --  0.7600141 -  0.7619619
     "11011011101110111011011101110110",  --  0.7620247 -  0.7639725
     "11101110110111011101110110111011",  --  0.7640353 -  0.7659831
     "10110111011101101110111011101101",  --  0.7660460 -  0.7679937
     "11011101101110111011101101110111",  --  0.7680566 -  0.7700044
     "01101110111011101101110111011101",  --  0.7700672 -  0.7720150
     "10111011101101110111011101101110",  --  0.7720778 -  0.7740256
     "11101110110111011101101110111011",  --  0.7740884 -  0.7760362
     "10110111011101110110111011101110",  --  0.7760990 -  0.7780468
     "11011101110111011011101110111011",  --  0.7781097 -  0.7800575
     "01110111011101101110111011101101",  --  0.7801203 -  0.7820681
     "11011101110110111011101110111011",  --  0.7821309 -  0.7840787
     "01110111011101101110111011101101",  --  0.7841415 -  0.7860893
     "11011101110111011011101110111011",  --  0.7861521 -  0.7880999
     "01110111011101110110111011101110",  --  0.7881628 -  0.7901106
     "11011101110111011101101110111011",  --  0.7901734 -  0.7921212
     "10111011011101110111011101101110",  --  0.7921840 -  0.7941318
     "11101110111011011101110111011101",  --  0.7941946 -  0.7961424
     "10111011101110111011011101110111",  --  0.7962052 -  0.7981530
     "01110110111011101110111011101101",  --  0.7982159 -  0.8001636
     "11011101110111011011101110111011",  --  0.8002265 -  0.8021743
     "10111011011101110111011101110110",  --  0.8022371 -  0.8041849
     "11101110111011101110110111011101",  --  0.8042477 -  0.8061955
     "11011101110110111011101110111011",  --  0.8062583 -  0.8082061
     "10111011011101110111011101110111",  --  0.8082690 -  0.8102167
     "01101110111011101110111011101101",  --  0.8102796 -  0.8122274
     "11011101110111011101110110111011",  --  0.8122902 -  0.8142380
     "10111011101110111011101101110111",  --  0.8143008 -  0.8162486
     "01110111011101110111011011101110",  --  0.8163114 -  0.8182592
     "11101110111011101110110111011101",  --  0.8183221 -  0.8202698
     "11011101110111011101110110111011",  --  0.8203327 -  0.8222805
     "10111011101110111011101110111011",  --  0.8223433 -  0.8242911
     "01110111011101110111011101110111",  --  0.8243539 -  0.8263017
     "01110110111011101110111011101110",  --  0.8263645 -  0.8283123
     "11101110111011101110110111011101",  --  0.8283752 -  0.8303229
     "11011101110111011101110111011101",  --  0.8303858 -  0.8323336
     "11011101110110111011101110111011",  --  0.8323964 -  0.8343442
     "10111011101110111011101110111011",  --  0.8344070 -  0.8363548
     "10111011101101110111011101110111",  --  0.8364176 -  0.8383654
     "01110111011101110111011101110111",  --  0.8384282 -  0.8403760
     "01110111011101110111011101110111",  --  0.8404389 -  0.8423867
     "01110110111011101110111011101110",  --  0.8424495 -  0.8443973
     "11101110111011101110111011101110",  --  0.8444601 -  0.8464079
     "11101110111011101110111011101110",  --  0.8464707 -  0.8484185
     "11101110111011101110111011101110",  --  0.8484813 -  0.8504291
     "11101110111011101110111011101110",  --  0.8504920 -  0.8524398
     "11101110111011101110111011101110",  --  0.8525026 -  0.8544504
     "11101110111011101110111011101110",  --  0.8545132 -  0.8564610
     "11101110111011101110111011101110",  --  0.8565238 -  0.8584716
     "11101110111011101110111011101110",  --  0.8585344 -  0.8604822
     "11101110111011101110111011101110",  --  0.8605451 -  0.8624928
     "11110111011101110111011101110111",  --  0.8625557 -  0.8645035
     "01110111011101110111011101110111",  --  0.8645663 -  0.8665141
     "01110111011101110111011101111011",  --  0.8665769 -  0.8685247
     "10111011101110111011101110111011",  --  0.8685875 -  0.8705353
     "10111011101110111011101110111101",  --  0.8705982 -  0.8725459
     "11011101110111011101110111011101",  --  0.8726088 -  0.8745566
     "11011101110111011110111011101110",  --  0.8746194 -  0.8765672
     "11101110111011101110111011101110",  --  0.8766300 -  0.8785778
     "11110111011101110111011101110111",  --  0.8786406 -  0.8805884
     "01110111011110111011101110111011",  --  0.8806513 -  0.8825990
     "10111011101110111011110111011101",  --  0.8826619 -  0.8846097
     "11011101110111011101110111101110",  --  0.8846725 -  0.8866203
     "11101110111011101110111011110111",  --  0.8866831 -  0.8886309
     "01110111011101110111011101111011",  --  0.8886937 -  0.8906415
     "10111011101110111011101111011101",  --  0.8907043 -  0.8926521
     "11011101110111011101111011101110",  --  0.8927150 -  0.8946628
     "11101110111011101111011101110111",  --  0.8947256 -  0.8966734
     "01110111011110111011101110111011",  --  0.8967362 -  0.8986840
     "10111101110111011101110111011110",  --  0.8987468 -  0.9006946
     "11101110111011101110111101110111",  --  0.9007574 -  0.9027052
     "01110111011101111011101110111011",  --  0.9027681 -  0.9047159
     "10111101110111011101110111101110",  --  0.9047787 -  0.9067265
     "11101110111011101111011101110111",  --  0.9067893 -  0.9087371
     "01110111101110111011101110111101",  --  0.9087999 -  0.9107477
     "11011101110111101110111011101110",  --  0.9108105 -  0.9127583
     "11110111011101110111011110111011",  --  0.9128212 -  0.9147689
     "10111011110111011101110111011110",  --  0.9148318 -  0.9167796
     "11101110111011110111011101110111",  --  0.9168424 -  0.9187902
     "10111011101110111011110111011101",  --  0.9188530 -  0.9208008
     "11011110111011101110111101110111",  --  0.9208636 -  0.9228114
     "01110111101110111011101111011101",  --  0.9228743 -  0.9248220
     "11011101111011101110111101110111",  --  0.9248849 -  0.9268327
     "01110111101110111011101111011101",  --  0.9268955 -  0.9288433
     "11011101111011101110111101110111",  --  0.9289061 -  0.9308539
     "01110111101110111011110111011101",  --  0.9309167 -  0.9328645
     "11011110111011101111011101110111",  --  0.9329274 -  0.9348751
     "01111011101110111101110111011101",  --  0.9349380 -  0.9368858
     "11101110111011110111011101111011",  --  0.9369486 -  0.9388964
     "10111011110111011101110111101110",  --  0.9389592 -  0.9409070
     "11101111011101110111101110111011",  --  0.9409698 -  0.9429176
     "11011101110111101110111011110111",  --  0.9429805 -  0.9449282
     "01110111101110111011110111011101",  --  0.9449911 -  0.9469389
     "11101110111011110111011101111011",  --  0.9470017 -  0.9489495
     "10111011110111011101111011101110",  --  0.9490123 -  0.9509601
     "11110111011110111011101111011101",  --  0.9510229 -  0.9529707
     "11011110111011101111011101110111",  --  0.9530335 -  0.9549813
     "10111011110111011101111011101110",  --  0.9550442 -  0.9569920
     "11110111011110111011101111011101",  --  0.9570548 -  0.9590026
     "11011110111011110111011101111011",  --  0.9590654 -  0.9610132
     "10111101110111011110111011110111",  --  0.9610760 -  0.9630238
     "01110111101110111101110111011110",  --  0.9630866 -  0.9650344
     "11101111011101110111101110111101",  --  0.9650973 -  0.9670451
     "11011101111011101111011101110111",  --  0.9671079 -  0.9690557
     "10111011110111011110111011101111",  --  0.9691185 -  0.9710663
     "01110111101110111101110111011110",  --  0.9711291 -  0.9730769
     "11101111011101111011101110111101",  --  0.9731397 -  0.9750875
     "11011110111011110111011110111011",  --  0.9751504 -  0.9770981
     "10111101110111101110111101110111",  --  0.9771610 -  0.9791088
     "10111011110111011101111011101111",  --  0.9791716 -  0.9811194
     "01110111101110111101110111101110",  --  0.9811822 -  0.9831300
     "11110111011110111011110111011101",  --  0.9831928 -  0.9851406
     "11101110111101110111101110111101",  --  0.9852035 -  0.9871512
     "11011110111011110111011110111011",  --  0.9872141 -  0.9891619
     "11011101111011101111011101111011",  --  0.9892247 -  0.9911725
     "10111101110111101110111101110111",  --  0.9912353 -  0.9931831
     "10111011110111011110111011110111",  --  0.9932459 -  0.9951937
     "01111011101111011101111011101111",  --  0.9952566 -  0.9972043
     "01110111101111011101111011101111",  --  0.9972672 -  0.9992150
     "01110111101110111101110111101110",  --  0.9992778 -  1.0012256
     "11110111011110111101110111101110",  --  1.0012884 -  1.0032362
     "11110111011110111011110111011110",  --  1.0032990 -  1.0052468
     "11110111011110111011110111011110",  --  1.0053096 -  1.0072574
     "11101111011110111011110111011110",  --  1.0073203 -  1.0092681
     "11101111011110111011110111011110",  --  1.0093309 -  1.0112787
     "11101111011110111011110111011110",  --  1.0113415 -  1.0132893
     "11101111011110111011110111011110",  --  1.0133521 -  1.0152999
     "11110111011110111011110111011110",  --  1.0153627 -  1.0173105
     "11110111011110111011110111101110",  --  1.0173734 -  1.0193212
     "11110111011110111101110111101111",  --  1.0193840 -  1.0213318
     "01110111101110111101111011101111",  --  1.0213946 -  1.0233424
     "01110111101111011101111011110111",  --  1.0234052 -  1.0253530
     "01111011101111011110111011110111",  --  1.0254158 -  1.0273636
     "10111011110111101110111101110111",  --  1.0274265 -  1.0293742
     "10111101110111101111011101111011",  --  1.0294371 -  1.0313849
     "11011101111011110111011110111011",  --  1.0314477 -  1.0333955
     "11011110111011110111101110111101",  --  1.0334583 -  1.0354061
     "11101110111101111011101111011110",  --  1.0354689 -  1.0374167
     "11101111011110111011110111101110",  --  1.0374796 -  1.0394273
     "11110111101111011101111011110111",  --  1.0394902 -  1.0414380
     "01111011110111011110111101110111",  --  1.0415008 -  1.0434486
     "10111101110111101111011110111011",  --  1.0435114 -  1.0454592
     "11011110111011110111101110111101",  --  1.0455220 -  1.0474698
     "11101111011101111011110111011110",  --  1.0475327 -  1.0494804
     "11110111101110111101111011101111",  --  1.0495433 -  1.0514911
     "01111011110111011110111101111011",  --  1.0515539 -  1.0535017
     "10111101111011101111011110111101",  --  1.0535645 -  1.0555123
     "11011110111101111011101111011110",  --  1.0555751 -  1.0575229
     "11110111011110111101111011101111",  --  1.0575858 -  1.0595335
     "01111011110111011110111101111011",  --  1.0595964 -  1.0615442
     "10111101111011110111011110111101",  --  1.0616070 -  1.0635548
     "11101110111101111011110111101110",  --  1.0636176 -  1.0655654
     "11110111101111011101111011110111",  --  1.0656282 -  1.0675760
     "10111101110111101111011110111011",  --  1.0676388 -  1.0695866
     "11011110111101111011101111011110",  --  1.0696495 -  1.0715973
     "11110111101110111101111011110111",  --  1.0716601 -  1.0736079
     "10111011110111101111011110111011",  --  1.0736707 -  1.0756185
     "11011110111101111011110111011110",  --  1.0756813 -  1.0776291
     "11110111101111011101111011110111",  --  1.0776919 -  1.0796397
     "10111101111011101111011110111101",  --  1.0797026 -  1.0816504
     "11101111011101111011110111101111",  --  1.0817132 -  1.0836610
     "01111011101111011110111101111011",  --  1.0837238 -  1.0856716
     "11011101111011110111101111011110",  --  1.0857344 -  1.0876822
     "11110111011110111101111011110111",  --  1.0877450 -  1.0896928
     "10111101110111101111011110111101",  --  1.0897557 -  1.0917034
     "11101111011110111011110111101111",  --  1.0917663 -  1.0937141
     "01111011110111101111011101111011",  --  1.0937769 -  1.0957247
     "11011110111101111011110111101111",  --  1.0957875 -  1.0977353
     "01110111101111011110111101111011",  --  1.0977981 -  1.0997459
     "11011110111101111011101111011110",  --  1.0998088 -  1.1017565
     "11110111101111011110111101111011",  --  1.1018194 -  1.1037672
     "11011110111011110111101111011110",  --  1.1038300 -  1.1057778
     "11110111101111011110111101111011",  --  1.1058406 -  1.1077884
     "11011101111011110111101111011110",  --  1.1078512 -  1.1097990
     "11110111101111011110111101111011",  --  1.1098619 -  1.1118096
     "11011110111101111011101111011110",  --  1.1118725 -  1.1138203
     "11110111101111011110111101111011",  --  1.1138831 -  1.1158309
     "11011110111101111011110111101111",  --  1.1158937 -  1.1178415
     "01111011110111101111011110111101",  --  1.1179043 -  1.1198521
     "11101111011110111101110111101111",  --  1.1199149 -  1.1218627
     "01111011110111101111011110111101",  --  1.1219256 -  1.1238734
     "11101111011110111101111011110111",  --  1.1239362 -  1.1258840
     "10111101111011110111101111011110",  --  1.1259468 -  1.1278946
     "11110111101111011110111101111011",  --  1.1279574 -  1.1299052
     "11011110111101111011110111101111",  --  1.1299680 -  1.1319158
     "01111011110111101111011110111101",  --  1.1319787 -  1.1339265
     "11101111011110111101111101111011",  --  1.1339893 -  1.1359371
     "11011110111101111011110111101111",  --  1.1359999 -  1.1379477
     "01111011110111101111011110111101",  --  1.1380105 -  1.1399583
     "11101111011110111101111011110111",  --  1.1400211 -  1.1419689
     "10111101111011110111110111101111",  --  1.1420318 -  1.1439795
     "01111011110111101111011110111101",  --  1.1440424 -  1.1459902
     "11101111011110111101111011110111",  --  1.1460530 -  1.1480008
     "10111110111101111011110111101111",  --  1.1480636 -  1.1500114
     "01111011110111101111011110111101",  --  1.1500742 -  1.1520220
     "11101111101111011110111101111011",  --  1.1520849 -  1.1540326
     "11011110111101111011110111101111",  --  1.1540955 -  1.1560433
     "10111101111011110111101111011110",  --  1.1561061 -  1.1580539
     "11110111101111011111011110111101",  --  1.1581167 -  1.1600645
     "11101111011110111101111011111011",  --  1.1601273 -  1.1620751
     "11011110111101111011110111101111",  --  1.1621380 -  1.1640857
     "01111011111011110111101111011110",  --  1.1641486 -  1.1660964
     "11110111101111101111011110111101",  --  1.1661592 -  1.1681070
     "11101111011110111110111101111011",  --  1.1681698 -  1.1701176
     "11011110111101111011111011110111",  --  1.1701804 -  1.1721282
     "10111101111011110111101111101111",  --  1.1721911 -  1.1741388
     "01111011110111101111011111011110",  --  1.1742017 -  1.1761495
     "11110111101111011110111110111101",  --  1.1762123 -  1.1781601
     "11101111011110111110111101111011",  --  1.1782229 -  1.1801707
     "11011110111101111101111011110111",  --  1.1802335 -  1.1821813
     "10111101111101111011110111101111",  --  1.1822441 -  1.1841919
     "01111101111011110111101111011111",  --  1.1842548 -  1.1862026
     "01111011110111101111011111011110",  --  1.1862654 -  1.1882132
     "11110111101111011111011110111101",  --  1.1882760 -  1.1902238
     "11101111011111011110111101111011",  --  1.1902866 -  1.1922344
     "11101111011110111101111011111011",  --  1.1922972 -  1.1942450
     "11011110111101111101111011110111",  --  1.1943079 -  1.1962557
     "10111110111101111011110111101111",  --  1.1963185 -  1.1982663
     "10111101111011110111110111101111",  --  1.1983291 -  1.2002769
     "01111011111011110111101111011111",  --  1.2003397 -  1.2022875
     "01111011110111101111101111011110",  --  1.2023503 -  1.2042981
     "11111011110111101111011111011110",  --  1.2043610 -  1.2063087
     "11110111101111101111011110111101",  --  1.2063716 -  1.2083194
     "11110111101111011111011110111101",  --  1.2083822 -  1.2103300
     "11101111101111011110111110111101",  --  1.2103928 -  1.2123406
     "11101111011111011110111101111101",  --  1.2124034 -  1.2143512
     "11101111011110111110111101111011",  --  1.2144141 -  1.2163618
     "11101111011110111110111101111011",  --  1.2164247 -  1.2183725
     "11101111011110111101111101111011",  --  1.2184353 -  1.2203831
     "11011111011110111101111101111011",  --  1.2204459 -  1.2223937
     "11011111011110111101111101111011",  --  1.2224565 -  1.2244043
     "11011111011110111101111101111011",  --  1.2244672 -  1.2264149
     "11011111011110111101111101111011",  --  1.2264778 -  1.2284256
     "11011111011110111101111101111011",  --  1.2284884 -  1.2304362
     "11011111011110111101111101111011",  --  1.2304990 -  1.2324468
     "11011111011110111101111101111011",  --  1.2325096 -  1.2344574
     "11101111011110111110111101111011",  --  1.2345202 -  1.2364680
     "11101111011110111110111101111101",  --  1.2365309 -  1.2384787
     "11101111011111011110111101111101",  --  1.2385415 -  1.2404893
     "11101111101111011110111110111101",  --  1.2405521 -  1.2424999
     "11101111101111011111011110111101",  --  1.2425627 -  1.2445105
     "11110111101111101111011110111110",  --  1.2445733 -  1.2465211
     "11110111110111101111011111011110",  --  1.2465840 -  1.2485318
     "11111011110111101111101111011111",  --  1.2485946 -  1.2505424
     "01111011110111110111101111101111",  --  1.2506052 -  1.2525530
     "01111011111011110111110111101111",  --  1.2526158 -  1.2545636
     "10111101111011111011110111110111",  --  1.2546264 -  1.2565742
     "10111110111101111011111011110111",  --  1.2566371 -  1.2585848
     "11011110111110111101111011111011",  --  1.2586477 -  1.2605955
     "11011111011110111110111101111101",  --  1.2606583 -  1.2626061
     "11101111011111011110111110111101",  --  1.2626689 -  1.2646167
     "11110111101111101111011111011110",  --  1.2646795 -  1.2666273
     "11110111110111101111101111011111",  --  1.2666902 -  1.2686379
     "01111011111011110111110111101111",  --  1.2687008 -  1.2706486
     "10111101111011111011110111110111",  --  1.2707114 -  1.2726592
     "10111110111101111101111011111011",  --  1.2727220 -  1.2746698
     "11011111011110111110111101111101",  --  1.2747326 -  1.2766804
     "11101111101111011111011110111110",  --  1.2767433 -  1.2786910
     "11110111110111101111101111011111",  --  1.2787539 -  1.2807017
     "01111011111011110111110111101111",  --  1.2807645 -  1.2827123
     "10111101111101111011111011110111",  --  1.2827751 -  1.2847229
     "11011110111110111101111101111011",  --  1.2847857 -  1.2867335
     "11101111011111011110111110111101",  --  1.2867964 -  1.2887441
     "11110111101111101111011111011110",  --  1.2888070 -  1.2907548
     "11111011110111110111110111101111",  --  1.2908176 -  1.2927654
     "10111101111101111011111011110111",  --  1.2928282 -  1.2947760
     "11011110111110111101111101111101",  --  1.2948388 -  1.2967866
     "11101111101111011111011110111110",  --  1.2968494 -  1.2987972
     "11110111110111101111101111101111",  --  1.2988601 -  1.3008079
     "01111101111011111011110111110111",  --  1.3008707 -  1.3028185
     "10111110111110111101111101111011",  --  1.3028813 -  1.3048291
     "11101111011111011111011110111110",  --  1.3048919 -  1.3068397
     "11110111110111101111101111101111",  --  1.3069025 -  1.3088503
     "01111101111011111011110111110111",  --  1.3089132 -  1.3108610
     "11011110111110111101111101111101",  --  1.3109238 -  1.3128716
     "11101111101111011111011110111110",  --  1.3129344 -  1.3148822
     "11111011110111110111101111101111",  --  1.3149450 -  1.3168928
     "10111101111101111011111011111011",  --  1.3169556 -  1.3189034
     "11011111011110111110111110111101",  --  1.3189663 -  1.3209140
     "11110111101111101111101111011111",  --  1.3209769 -  1.3229247
     "01111101111011111011110111110111",  --  1.3229875 -  1.3249353
     "11011110111110111101111101111101",  --  1.3249981 -  1.3269459
     "11101111101111101111011111011110",  --  1.3270087 -  1.3289565
     "11111011111011110111110111110111",  --  1.3290194 -  1.3309671
     "10111110111110111101111101111011",  --  1.3310300 -  1.3329778
     "11101111101111011111011111011110",  --  1.3330406 -  1.3349884
     "11111011111011110111110111110111",  --  1.3350512 -  1.3369990
     "10111110111101111101111101111011",  --  1.3370618 -  1.3390096
     "11101111101111011111011111011110",  --  1.3390725 -  1.3410202
     "11111011111011110111110111110111",  --  1.3410831 -  1.3430309
     "10111110111110111101111101111101",  --  1.3430937 -  1.3450415
     "11101111101111101111011111011111",  --  1.3451043 -  1.3470521
     "01111011111011111011110111110111",  --  1.3471149 -  1.3490627
     "11011110111110111110111101111101",  --  1.3491255 -  1.3510733
     "11110111110111101111101111101111",  --  1.3511362 -  1.3530840
     "01111101111101111011111011111011",  --  1.3531468 -  1.3550946
     "11011111011111011110111110111110",  --  1.3551574 -  1.3571052
     "11111011110111110111110111101111",  --  1.3571680 -  1.3591158
     "10111110111101111101111101111101",  --  1.3591786 -  1.3611264
     "11101111101111101111011111011111",  --  1.3611893 -  1.3631371
     "01111101111011111011111011110111",  --  1.3631999 -  1.3651477
     "11011111011111011110111110111110",  --  1.3652105 -  1.3671583
     "11110111110111110111110111101111",  --  1.3672211 -  1.3691689
     "10111110111101111101111101111101",  --  1.3692317 -  1.3711795
     "11101111101111101111101111011111",  --  1.3712424 -  1.3731901
     "01111101111011111011111011111011",  --  1.3732530 -  1.3752008
     "11011111011111011111011110111110",  --  1.3752636 -  1.3772114
     "11111011111011110111110111110111",  --  1.3772742 -  1.3792220
     "11011110111110111110111110111101",  --  1.3792848 -  1.3812326
     "11110111110111110111101111101111",  --  1.3812955 -  1.3832432
     "10111110111101111101111101111101",  --  1.3833061 -  1.3852539
     "11101111101111101111101111011111",  --  1.3853167 -  1.3872645
     "01111101111101111011111011111011",  --  1.3873273 -  1.3892751
     "11101111011111011111011111011111",  --  1.3893379 -  1.3912857
     "01111011111011111011111011110111",  --  1.3913486 -  1.3932963
     "11011111011111011110111110111110",  --  1.3933592 -  1.3953070
     "11111011111011110111110111110111",  --  1.3953698 -  1.3973176
     "11011110111110111110111110111110",  --  1.3973804 -  1.3993282
     "11110111110111110111110111110111",  --  1.3993910 -  1.4013388
     "10111110111110111110111110111101",  --  1.4014017 -  1.4033494
     "11110111110111110111101111101111",  --  1.4034123 -  1.4053601
     "10111110111110111101111101111101",  --  1.4054229 -  1.4073707
     "11110111110111101111101111101111",  --  1.4074335 -  1.4093813
     "10111110111101111101111101111101",  --  1.4094441 -  1.4113919
     "11110111110111101111101111101111",  --  1.4114547 -  1.4134025
     "10111110111101111101111101111101",  --  1.4134654 -  1.4154132
     "11110111101111101111101111101111",  --  1.4154760 -  1.4174238
     "10111110111101111101111101111101",  --  1.4174866 -  1.4194344
     "11110111101111101111101111101111",  --  1.4194972 -  1.4214450
     "10111110111101111101111101111101",  --  1.4215078 -  1.4234556
     "11110111110111101111101111101111",  --  1.4235185 -  1.4254663
     "10111110111101111101111101111101",  --  1.4255291 -  1.4274769
     "11110111110111110111101111101111",  --  1.4275397 -  1.4294875
     "10111110111110111110111101111101",  --  1.4295503 -  1.4314981
     "11110111110111110111110111101111",  --  1.4315609 -  1.4335087
     "10111110111110111110111110111101",  --  1.4335716 -  1.4355193
     "11110111110111110111110111110111",  --  1.4355822 -  1.4375300
     "11011110111110111110111110111110",  --  1.4375928 -  1.4395406
     "11111011111011110111110111110111",  --  1.4396034 -  1.4415512
     "11011111011111011111011110111110",  --  1.4416140 -  1.4435618
     "11111011111011111011111011111011",  --  1.4436247 -  1.4455724
     "11011111011111011111011111011111",  --  1.4456353 -  1.4475831
     "01111101111011111011111011111011",  --  1.4476459 -  1.4495937
     "11101111101111101111101111011111",  --  1.4496565 -  1.4516043
     "01111101111101111101111101111101",  --  1.4516671 -  1.4536149
     "11101111101111101111101111101111",  --  1.4536778 -  1.4556255
     "10111110111110111101111101111101",  --  1.4556884 -  1.4576362
     "11110111110111110111110111110111",  --  1.4576990 -  1.4596468
     "11011110111110111110111110111110",  --  1.4597096 -  1.4616574
     "11111011111011111011110111110111",  --  1.4617202 -  1.4636680
     "11011111011111011111011111011111",  --  1.4637308 -  1.4656786
     "01111101111011111011111011111011",  --  1.4657415 -  1.4676893
     "11101111101111101111101111101111",  --  1.4677521 -  1.4696999
     "01111101111101111101111101111101",  --  1.4697627 -  1.4717105
     "11110111110111110111110111101111",  --  1.4717733 -  1.4737211
     "10111110111110111110111110111110",  --  1.4737839 -  1.4757317
     "11111011111011111011110111110111",  --  1.4757946 -  1.4777424
     "11011111011111011111011111011111",  --  1.4778052 -  1.4797530
     "01111101111101111011111011111011",  --  1.4798158 -  1.4817636
     "11101111101111101111101111101111",  --  1.4818264 -  1.4837742
     "10111110111110111101111101111101",  --  1.4838370 -  1.4857848
     "11110111110111110111110111110111",  --  1.4858477 -  1.4877954
     "11011111011111011110111110111110",  --  1.4878583 -  1.4898061
     "11111011111011111011111011111011",  --  1.4898689 -  1.4918167
     "11101111101111101111101111011111",  --  1.4918795 -  1.4938273
     "01111101111101111101111101111101",  --  1.4938901 -  1.4958379
     "11110111110111110111110111110111",  --  1.4959008 -  1.4978485
     "10111110111110111110111110111110",  --  1.4979114 -  1.4998592
     "11111011111011111011111011111011",  --  1.4999220 -  1.5018698
     "11101111101111011111011111011111",  --  1.5019326 -  1.5038804
     "01111101111101111101111101111101",  --  1.5039432 -  1.5058910
     "11110111110111110111110111110111",  --  1.5059539 -  1.5079016
     "10111110111110111110111110111110",  --  1.5079645 -  1.5099123
     "11111011111011111011111011111011",  --  1.5099751 -  1.5119229
     "11101111101111101111101111011111",  --  1.5119857 -  1.5139335
     "01111101111101111101111101111101",  --  1.5139963 -  1.5159441
     "11110111110111110111110111110111",  --  1.5160070 -  1.5179547
     "11011111011111011110111110111110",  --  1.5180176 -  1.5199654
     "11111011111011111011111011111011",  --  1.5200282 -  1.5219760
     "11101111101111101111101111101111",  --  1.5220388 -  1.5239866
     "10111110111110111101111101111101",  --  1.5240494 -  1.5259972
     "11110111110111110111110111110111",  --  1.5260600 -  1.5280078
     "11011111011111011111011111011111",  --  1.5280707 -  1.5300185
     "01111101111101111101111011111011",  --  1.5300813 -  1.5320291
     "11101111101111101111101111101111",  --  1.5320919 -  1.5340397
     "10111110111110111110111110111110",  --  1.5341025 -  1.5360503
     "11111011111011111011111011111011",  --  1.5361131 -  1.5380609
     "11011111011111011111011111011111",  --  1.5381238 -  1.5400716
     "01111101111101111101111101111101",  --  1.5401344 -  1.5420822
     "11110111110111110111110111110111",  --  1.5421450 -  1.5440928
     "11011111011111011110111110111110",  --  1.5441556 -  1.5461034
     "11111011111011111011111011111011",  --  1.5461662 -  1.5481140
     "11101111101111101111101111101111",  --  1.5481769 -  1.5501246
     "10111110111110111110111110111110",  --  1.5501875 -  1.5521353
     "11111011110111110111110111110111",  --  1.5521981 -  1.5541459
     "11011111011111011111011111011111",  --  1.5542087 -  1.5561565
     "01111101111101111101111101111101",  --  1.5562193 -  1.5581671
     "11110111110111110111110111110111",  --  1.5582300 -  1.5601777
     "11011110111110111110111110111110",  --  1.5602406 -  1.5621884
     "11111011111011111011111011111011",  --  1.5622512 -  1.5641990
     "11101111101111101111101111101111",  --  1.5642618 -  1.5662096
     "10111110111110111110111110111110",  --  1.5662724 -  1.5682202
     "11110111110111110111110111110111",  --  1.5682831 -  1.5702308
     "11011111011111011111011111011111",  --  1.5702937 -  1.5722415
     "01111101111101111101111101111101",  --  1.5723043 -  1.5742521
     "11110111110111110111110111101111",  --  1.5743149 -  1.5762627
     "10111110111110111110111110111110",  --  1.5763255 -  1.5782733
     "11111011111011111011111011111011",  --  1.5783361 -  1.5802839
     "11101111101111101111101111101111",  --  1.5803468 -  1.5822946
     "10111110111110111110111101111101",  --  1.5823574 -  1.5843052
     "11110111110111110111110111110111",  --  1.5843680 -  1.5863158
     "11011111011111011111011111011111",  --  1.5863786 -  1.5883264
     "01111101111101111101111101111101",  --  1.5883892 -  1.5903370
     "11110111110111110111101111101111",  --  1.5903999 -  1.5923477
     "10111110111110111110111110111110",  --  1.5924105 -  1.5943583
     "11111011111011111011111011111011",  --  1.5944211 -  1.5963689
     "11101111101111101111101111101111",  --  1.5964317 -  1.5983795
     "10111101111101111101111101111101",  --  1.5984423 -  1.6003901
     "11110111110111110111110111110111",  --  1.6004530 -  1.6024007
     "11011111011111011111011111011111",  --  1.6024636 -  1.6044114
     "01111101111101111101111011111011",  --  1.6044742 -  1.6064220
     "11101111101111101111101111101111",  --  1.6064848 -  1.6084326
     "10111110111110111110111110111110",  --  1.6084954 -  1.6104432
     "11111011111011111011111011111011",  --  1.6105061 -  1.6124538
     "11011111011111011111011111011111",  --  1.6125167 -  1.6144645
     "01111101111101111101111101111101",  --  1.6145273 -  1.6164751
     "11110111110111110111110111110111",  --  1.6165379 -  1.6184857
     "10111110111110111110111110111110",  --  1.6185485 -  1.6204963
     "11111011111011111011111011111011",  --  1.6205592 -  1.6225069
     "11101111101111101111101111101111",  --  1.6225698 -  1.6245176
     "01111101111101111101111101111101",  --  1.6245804 -  1.6265282
     "11110111110111110111110111110111",  --  1.6265910 -  1.6285388
     "11011111011111011111011110111110",  --  1.6286016 -  1.6305494
     "11111011111011111011111011111011",  --  1.6306123 -  1.6325600
     "11101111101111101111101111101111",  --  1.6326229 -  1.6345707
     "10111110111110111101111101111101",  --  1.6346335 -  1.6365813
     "11110111110111110111110111110111",  --  1.6366441 -  1.6385919
     "11011111011111011111011111011110",  --  1.6386547 -  1.6406025
     "11111011111011111011111011111011",  --  1.6406653 -  1.6426131
     "11101111101111101111101111101111",  --  1.6426760 -  1.6446238
     "10111110111101111101111101111101",  --  1.6446866 -  1.6466344
     "11110111110111110111110111110111",  --  1.6466972 -  1.6486450
     "11011111011111011110111110111110",  --  1.6487078 -  1.6506556
     "11111011111011111011111011111011",  --  1.6507184 -  1.6526662
     "11101111101111101111101111011111",  --  1.6527291 -  1.6546769
     "01111101111101111101111101111101",  --  1.6547397 -  1.6566875
     "11110111110111110111110111101111",  --  1.6567503 -  1.6586981
     "10111110111110111110111110111110",  --  1.6587609 -  1.6607087
     "11111011111011111011111011110111",  --  1.6607715 -  1.6627193
     "11011111011111011111011111011111",  --  1.6627822 -  1.6647299
     "01111101111101111101111011111011",  --  1.6647928 -  1.6667406
     "11101111101111101111101111101111",  --  1.6668034 -  1.6687512
     "10111110111101111101111101111101",  --  1.6688140 -  1.6707618
     "11110111110111110111110111110111",  --  1.6708246 -  1.6727724
     "11011110111110111110111110111110",  --  1.6728353 -  1.6747830
     "11111011111011111011111011110111",  --  1.6748459 -  1.6767937
     "11011111011111011111011111011111",  --  1.6768565 -  1.6788043
     "01111101111101111011111011111011",  --  1.6788671 -  1.6808149
     "11101111101111101111101111101111",  --  1.6808777 -  1.6828255
     "01111101111101111101111101111101",  --  1.6828884 -  1.6848361
     "11110111110111101111101111101111",  --  1.6848990 -  1.6868468
     "10111110111110111110111110111101",  --  1.6869096 -  1.6888574
     "11110111110111110111110111110111",  --  1.6889202 -  1.6908680
     "11011111011110111110111110111110",  --  1.6909308 -  1.6928786
     "11111011111011111011110111110111",  --  1.6929414 -  1.6948892
     "11011111011111011111011111011111",  --  1.6949521 -  1.6968999
     "01111011111011111011111011111011",  --  1.6969627 -  1.6989105
     "11101111101111011111011111011111",  --  1.6989733 -  1.7009211
     "01111101111101111101111011111011",  --  1.7009839 -  1.7029317
     "11101111101111101111101111011111",  --  1.7029945 -  1.7049423
     "01111101111101111101111101111101",  --  1.7050052 -  1.7069530
     "11101111101111101111101111101111",  --  1.7070158 -  1.7089636
     "10111101111101111101111101111101",  --  1.7090264 -  1.7109742
     "11110111101111101111101111101111",  --  1.7110370 -  1.7129848
     "10111110111110111101111101111101",  --  1.7130476 -  1.7149954
     "11110111110111110111101111101111",  --  1.7150583 -  1.7170060
     "10111110111110111101111101111101",  --  1.7170689 -  1.7190167
     "11110111110111110111101111101111",  --  1.7190795 -  1.7210273
     "10111110111110111110111101111101",  --  1.7210901 -  1.7230379
     "11110111110111110111101111101111",  --  1.7231007 -  1.7250485
     "10111110111110111110111101111101",  --  1.7251114 -  1.7270591
     "11110111110111110111101111101111",  --  1.7271220 -  1.7290698
     "10111110111110111101111101111101",  --  1.7291326 -  1.7310804
     "11110111110111101111101111101111",  --  1.7311432 -  1.7330910
     "10111110111101111101111101111101",  --  1.7331538 -  1.7351016
     "11110111101111101111101111101111",  --  1.7351645 -  1.7371122
     "10111101111101111101111101111101",  --  1.7371751 -  1.7391229
     "11101111101111101111101111101111",  --  1.7391857 -  1.7411335
     "01111101111101111101111101111011",  --  1.7411963 -  1.7431441
     "11101111101111101111011111011111",  --  1.7432069 -  1.7451547
     "01111101111101111011111011111011",  --  1.7452176 -  1.7471653
     "11101111011111011111011111011111",  --  1.7472282 -  1.7491760
     "01111011111011111011111011110111",  --  1.7492388 -  1.7511866
     "11011111011111011110111110111110",  --  1.7512494 -  1.7531972
     "11111011110111110111110111110111",  --  1.7532600 -  1.7552078
     "11011110111110111110111110111101",  --  1.7552706 -  1.7572184
     "11110111110111110111101111101111",  --  1.7572813 -  1.7592291
     "10111110111101111101111101111101",  --  1.7592919 -  1.7612397
     "11101111101111101111101111011111",  --  1.7613025 -  1.7632503
     "01111101111101111011111011111011",  --  1.7633131 -  1.7652609
     "11011111011111011111011110111110",  --  1.7653237 -  1.7672715
     "11111011111011110111110111110111",  --  1.7673344 -  1.7692822
     "11011110111110111110111101111101",  --  1.7693450 -  1.7712928
     "11110111110111101111101111101111",  --  1.7713556 -  1.7733034
     "10111101111101111101111011111011",  --  1.7733662 -  1.7753140
     "11101111101111011111011111011110",  --  1.7753768 -  1.7773246
     "11111011111011111011110111110111",  --  1.7773875 -  1.7793352
     "11011110111110111110111110111101",  --  1.7793981 -  1.7813459
     "11110111110111101111101111101111",  --  1.7814087 -  1.7833565
     "01111101111101111101111011111011",  --  1.7834193 -  1.7853671
     "11101111011111011111011110111110",  --  1.7854299 -  1.7873777
     "11111011110111110111110111101111",  --  1.7874406 -  1.7893883
     "10111110111110111101111101111101",  --  1.7894512 -  1.7913990
     "11101111101111101111011111011111",  --  1.7914618 -  1.7934096
     "01111011111011111011110111110111",  --  1.7934724 -  1.7954202
     "11011110111110111110111101111101",  --  1.7954830 -  1.7974308
     "11110111101111101111101111011111",  --  1.7974937 -  1.7994414
     "01111101111011111011111011110111",  --  1.7995043 -  1.8014521
     "11011111011110111110111110111101",  --  1.8015149 -  1.8034627
     "11110111110111101111101111011111",  --  1.8035255 -  1.8054733
     "01111101111011111011111011110111",  --  1.8055361 -  1.8074839
     "11011111011110111110111110111101",  --  1.8075467 -  1.8094945
     "11110111101111101111101111011111",  --  1.8095574 -  1.8115052
     "01111101111011111011111011110111",  --  1.8115680 -  1.8135158
     "11011110111110111110111101111101",  --  1.8135786 -  1.8155264
     "11110111101111101111011111011111",  --  1.8155892 -  1.8175370
     "01111011111011110111110111110111",  --  1.8175998 -  1.8195476
     "10111110111110111101111101111011",  --  1.8196105 -  1.8215583
     "11101111101111011111011110111110",  --  1.8216211 -  1.8235689
     "11111011110111110111101111101111",  --  1.8236317 -  1.8255795
     "10111101111101111011111011111011",  --  1.8256423 -  1.8275901
     "11011111011110111110111101111101",  --  1.8276529 -  1.8296007
     "11110111101111101111011111011111",  --  1.8296636 -  1.8316113
     "01111011111011110111110111101111",  --  1.8316742 -  1.8336220
     "10111110111101111101111011111011",  --  1.8336848 -  1.8356326
     "11011111011111011110111110111101",  --  1.8356954 -  1.8376432
     "11110111101111101111011111011111",  --  1.8377060 -  1.8396538
     "01111011111011110111110111101111",  --  1.8397167 -  1.8416644
     "10111101111101111101111011111011",  --  1.8417273 -  1.8436751
     "11011111011110111110111101111101",  --  1.8437379 -  1.8456857
     "11101111101111101111011111011110",  --  1.8457485 -  1.8476963
     "11111011110111110111101111101111",  --  1.8477591 -  1.8497069
     "01111101111011111011110111110111",  --  1.8497698 -  1.8517175
     "11011110111110111101111101111011",  --  1.8517804 -  1.8537282
     "11101111011111011110111110111101",  --  1.8537910 -  1.8557388
     "11110111101111101111011111011110",  --  1.8558016 -  1.8577494
     "11111011110111110111101111101111",  --  1.8578122 -  1.8597600
     "01111101111011111011110111110111",  --  1.8598229 -  1.8617706
     "10111110111101111101111011111011",  --  1.8618335 -  1.8637813
     "11011111011110111110111101111101",  --  1.8638441 -  1.8657919
     "11101111101111011111011110111110",  --  1.8658547 -  1.8678025
     "11110111110111101111101111011110",  --  1.8678653 -  1.8698131
     "11111011110111110111101111101111",  --  1.8698759 -  1.8718237
     "01111101111011111011110111110111",  --  1.8718866 -  1.8738344
     "10111110111101111011111011110111",  --  1.8738972 -  1.8758450
     "11011110111110111101111101111011",  --  1.8759078 -  1.8778556
     "11101111011110111110111101111101",  --  1.8779184 -  1.8798662
     "11101111101111011110111110111101",  --  1.8799290 -  1.8818768
     "11110111101111101111011111011110",  --  1.8819397 -  1.8838875
     "11110111110111101111101111011111",  --  1.8839503 -  1.8858981
     "01111011110111110111101111101111",  --  1.8859609 -  1.8879087
     "01111011111011110111110111101111",  --  1.8879715 -  1.8899193
     "10111101111011111011110111110111",  --  1.8899821 -  1.8919299
     "10111101111101111011111011110111",  --  1.8919928 -  1.8939405
     "10111110111101111101111011110111",  --  1.8940034 -  1.8959512
     "11011110111110111101111011111011",  --  1.8960140 -  1.8979618
     "11011111011110111101111101111011",  --  1.8980246 -  1.8999724
     "11011111011110111110111101111011",  --  1.9000352 -  1.9019830
     "11101111011110111110111101111101",  --  1.9020459 -  1.9039936
     "11101111011111011110111101111101",  --  1.9040565 -  1.9060043
     "11101111011111011110111110111101",  --  1.9060671 -  1.9080149
     "11101111101111011110111110111101",  --  1.9080777 -  1.9100255
     "11101111101111011110111110111101",  --  1.9100883 -  1.9120361
     "11101111101111011110111110111101",  --  1.9120990 -  1.9140467
     "11110111101111011111011110111101",  --  1.9141096 -  1.9160574
     "11110111101111011110111110111101",  --  1.9161202 -  1.9180680
     "11101111101111011110111110111101",  --  1.9181308 -  1.9200786
     "11101111101111011110111110111101",  --  1.9201414 -  1.9220892
     "11101111101111011110111110111101",  --  1.9221520 -  1.9240998
     "11101111011111011110111101111101",  --  1.9241627 -  1.9261105
     "11101111011111011110111101111011",  --  1.9261733 -  1.9281211
     "11101111011110111110111101111011",  --  1.9281839 -  1.9301317
     "11011111011110111101111101111011",  --  1.9301945 -  1.9321423
     "11011110111110111101111011110111",  --  1.9322051 -  1.9341529
     "11011110111101111101111011110111",  --  1.9342158 -  1.9361636
     "10111110111101111011110111110111",  --  1.9362264 -  1.9381742
     "10111101111011111011110111101111",  --  1.9382370 -  1.9401848
     "01111101111011110111101111101111",  --  1.9402476 -  1.9421954
     "01111011110111110111101111011110",  --  1.9422582 -  1.9442060
     "11111011110111101111011111011110",  --  1.9442689 -  1.9462166
     "11110111101111101111011110111101",  --  1.9462795 -  1.9482273
     "11101111101111011110111101111101",  --  1.9482901 -  1.9502379
     "11101111011110111101111101111011",  --  1.9503007 -  1.9522485
     "11011110111101111101111011110111",  --  1.9523113 -  1.9542591
     "10111110111101111011110111101111",  --  1.9543220 -  1.9562697
     "10111101111011110111101111011111",  --  1.9563326 -  1.9582804
     "01111011110111101111011111011110",  --  1.9583432 -  1.9602910
     "11110111101111011111011110111101",  --  1.9603538 -  1.9623016
     "11101111011110111110111101111011",  --  1.9623644 -  1.9643122
     "11011110111101111101111011110111",  --  1.9643751 -  1.9663228
     "10111101111011111011110111101111",  --  1.9663857 -  1.9683335
     "01111011110111110111101111011110",  --  1.9683963 -  1.9703441
     "11110111101111011111011110111101",  --  1.9704069 -  1.9723547
     "11101111011110111101111101111011",  --  1.9724175 -  1.9743653
     "11011110111101111011110111110111",  --  1.9744282 -  1.9763759
     "10111101111011110111101111011110",  --  1.9764388 -  1.9783866
     "11111011110111101111011110111101",  --  1.9784494 -  1.9803972
     "11101111011110111110111101111011",  --  1.9804600 -  1.9824078
     "11011110111101111011110111101111",  --  1.9824706 -  1.9844184
     "10111101111011110111101111011110",  --  1.9844812 -  1.9864290
     "11110111101111011111011110111101",  --  1.9864919 -  1.9884397
     "11101111011110111101111011110111",  --  1.9885025 -  1.9904503
     "10111101111011111011110111101111",  --  1.9905131 -  1.9924609
     "01111011110111101111011110111101",  --  1.9925237 -  1.9944715
     "11101111011110111101111101111011",  --  1.9945343 -  1.9964821
     "11011110111101111011110111101111",  --  1.9965450 -  1.9984928
     "01111011110111101111011110111101",  --  1.9985556 -  2.0005034
     "11101111011110111101111011111011",  --  2.0005662 -  2.0025140
     "11011110111101111011110111101111",  --  2.0025768 -  2.0045246
     "01111011110111101111011110111101",  --  2.0045874 -  2.0065352
     "11101111011110111101111011110111",  --  2.0065981 -  2.0085458
     "10111101111011110111101111011110",  --  2.0086087 -  2.0105565
     "11110111101111011110111101111011",  --  2.0106193 -  2.0125671
     "11011110111101111011110111101111",  --  2.0126299 -  2.0145777
     "01111011110111101111011110111101",  --  2.0146405 -  2.0165883
     "11101111011110111101111011110111",  --  2.0166512 -  2.0185989
     "10111101111011110111101111011110",  --  2.0186618 -  2.0206096
     "11110111101111011110111101111011",  --  2.0206724 -  2.0226202
     "11011110111101111011110111101111",  --  2.0226830 -  2.0246308
     "01110111101111011110111101111011",  --  2.0246936 -  2.0266414
     "11011110111101111011110111101111",  --  2.0267043 -  2.0286520
     "01111011110111101111011110111101",  --  2.0287149 -  2.0306627
     "11011110111101111011110111101111",  --  2.0307255 -  2.0326733
     "01111011110111101111011110111101",  --  2.0327361 -  2.0346839
     "11101111011101111011110111101111",  --  2.0347467 -  2.0366945
     "01111011110111101111011110111101",  --  2.0367573 -  2.0387051
     "11101110111101111011110111101111",  --  2.0387680 -  2.0407158
     "01111011110111101111011101111011",  --  2.0407786 -  2.0427264
     "11011110111101111011110111101111",  --  2.0427892 -  2.0447370
     "01110111101111011110111101111011",  --  2.0447998 -  2.0467476
     "11011110111101110111101111011110",  --  2.0468104 -  2.0487582
     "11110111101111011101111011110111",  --  2.0488211 -  2.0507689
     "10111101111011110111101110111101",  --  2.0508317 -  2.0527795
     "11101111011110111101111011101111",  --  2.0528423 -  2.0547901
     "01111011110111101111011101111011",  --  2.0548529 -  2.0568007
     "11011110111101111011110111011110",  --  2.0568635 -  2.0588113
     "11110111101111011110111011110111",  --  2.0588742 -  2.0608219
     "10111101111011110111011110111101",  --  2.0608848 -  2.0628326
     "11101111011101111011110111101111",  --  2.0628954 -  2.0648432
     "01111011101111011110111101111011",  --  2.0649060 -  2.0668538
     "10111101111011110111101110111101",  --  2.0669166 -  2.0688644
     "11101111011110111011110111101111",  --  2.0689273 -  2.0708750
     "01111011101111011110111101111011",  --  2.0709379 -  2.0728857
     "10111101111011110111011110111101",  --  2.0729485 -  2.0748963
     "11101111011101111011110111101110",  --  2.0749591 -  2.0769069
     "11110111101111011110111011110111",  --  2.0769697 -  2.0789175
     "10111101110111101111011110111011",  --  2.0789804 -  2.0809281
     "11011110111101110111101111011110",  --  2.0809910 -  2.0829388
     "11101111011110111101110111101111",  --  2.0830016 -  2.0849494
     "01111011101111011110111101110111",  --  2.0850122 -  2.0869600
     "10111101110111101111011110111011",  --  2.0870228 -  2.0889706
     "11011110111101110111101111011101",  --  2.0890335 -  2.0909812
     "11101111011110111011110111101110",  --  2.0910441 -  2.0929919
     "11110111101111011101111011110111",  --  2.0930547 -  2.0950025
     "01111011110111101110111101111011",  --  2.0950653 -  2.0970131
     "10111101111011101111011110111011",  --  2.0970759 -  2.0990237
     "11011110111101110111101111011101",  --  2.0990865 -  2.1010343
     "11101111011101111011110111011110",  --  2.1010972 -  2.1030450
     "11110111011110111101110111101111",  --  2.1031078 -  2.1050556
     "01110111101111011101111011110111",  --  2.1051184 -  2.1070662
     "01111011110111011110111101110111",  --  2.1071290 -  2.1090768
     "10111101110111101111011101111011",  --  2.1091396 -  2.1110874
     "10111101111011101111011110111011",  --  2.1111503 -  2.1130981
     "11011110111011110111101110111101",  --  2.1131609 -  2.1151087
     "11011110111101110111101111011101",  --  2.1151715 -  2.1171193
     "11101110111101111011101111011101",  --  2.1171821 -  2.1191299
     "11101111011101111011110111011110",  --  2.1191927 -  2.1211405
     "11101111011110111011110111011110",  --  2.1212034 -  2.1231511
     "11110111011110111011110111101110",  --  2.1232140 -  2.1251618
     "11110111011110111101110111101110",  --  2.1252246 -  2.1271724
     "11110111011110111101110111101110",  --  2.1272352 -  2.1291830
     "11110111101110111101110111101110",  --  2.1292458 -  2.1311936
     "11110111101110111101110111101110",  --  2.1312565 -  2.1332042
     "11110111011110111101110111101110",  --  2.1332671 -  2.1352149
     "11110111011110111101110111101110",  --  2.1352777 -  2.1372255
     "11110111011110111011110111011110",  --  2.1372883 -  2.1392361
     "11110111011110111011110111011110",  --  2.1392989 -  2.1412467
     "11101111011101111011101111011101",  --  2.1413096 -  2.1432573
     "11101110111101111011101111011101",  --  2.1433202 -  2.1452680
     "11101110111101110111101110111101",  --  2.1453308 -  2.1472786
     "11011110111011110111011110111011",  --  2.1473414 -  2.1492892
     "11011101111011101111011101111011",  --  2.1493520 -  2.1512998
     "10111101110111101110111101110111",  --  2.1513626 -  2.1533104
     "10111011110111011110111011110111",  --  2.1533733 -  2.1553211
     "01111011101111011101111011101110",  --  2.1553839 -  2.1573317
     "11110111011110111011110111011110",  --  2.1573945 -  2.1593423
     "11101111011101111011101111011101",  --  2.1594051 -  2.1613529
     "11011110111011110111011110111011",  --  2.1614157 -  2.1633635
     "11011101111011101110111101110111",  --  2.1634264 -  2.1653742
     "10111011110111011110111011101111",  --  2.1654370 -  2.1673848
     "01110111101110111101110111011110",  --  2.1674476 -  2.1693954
     "11101111011101111011101110111101",  --  2.1694582 -  2.1714060
     "11011110111011110111011101111011",  --  2.1714688 -  2.1734166
     "10111101110111011110111011110111",  --  2.1734795 -  2.1754272
     "01111011101110111101110111101110",  --  2.1754901 -  2.1774379
     "11101111011101111011101110111101",  --  2.1775007 -  2.1794485
     "11011110111011101111011101110111",  --  2.1795113 -  2.1814591
     "10111011110111011101111011101111",  --  2.1815219 -  2.1834697
     "01110111011110111011101111011101",  --  2.1835326 -  2.1854803
     "11101110111011110111011101111011",  --  2.1855432 -  2.1874910
     "10111011110111011110111011101111",  --  2.1875538 -  2.1895016
     "01110111011110111011101111011101",  --  2.1895644 -  2.1915122
     "11011110111011101111011101111011",  --  2.1915750 -  2.1935228
     "10111011110111011101111011101110",  --  2.1935857 -  2.1955334
     "11110111011101111011101110111101",  --  2.1955963 -  2.1975441
     "11011101111011101110111011110111",  --  2.1976069 -  2.1995547
     "01110111101110111011110111011101",  --  2.1996175 -  2.2015653
     "11101110111011110111011101111011",  --  2.2016281 -  2.2035759
     "10111011101111011101110111101110",  --  2.2036388 -  2.2055865
     "11101111011101110111011110111011",  --  2.2056494 -  2.2075972
     "10111101110111011101111011101110",  --  2.2076600 -  2.2096078
     "11110111011101110111101110111011",  --  2.2096706 -  2.2116184
     "11011101110111011110111011101110",  --  2.2116812 -  2.2136290
     "11110111011101110111101110111011",  --  2.2136918 -  2.2156396
     "11011101110111011110111011101110",  --  2.2157025 -  2.2176503
     "11110111011101110111101110111011",  --  2.2177131 -  2.2196609
     "10111101110111011101111011101110",  --  2.2197237 -  2.2216715
     "11101111011101110111011101111011",  --  2.2217343 -  2.2236821
     "10111011101111011101110111011110",  --  2.2237449 -  2.2256927
     "11101110111011101111011101110111",  --  2.2257556 -  2.2277034
     "01111011101110111011101111011101",  --  2.2277662 -  2.2297140
     "11011101110111101110111011101110",  --  2.2297768 -  2.2317246
     "11110111011101110111011110111011",  --  2.2317874 -  2.2337352
     "10111011101111011101110111011101",  --  2.2337980 -  2.2357458
     "11101110111011101110111101110111",  --  2.2358087 -  2.2377564
     "01110111011101111011101110111011",  --  2.2378193 -  2.2397671
     "10111011110111011101110111011110",  --  2.2398299 -  2.2417777
     "11101110111011101110111011110111",  --  2.2418405 -  2.2437883
     "01110111011101110111101110111011",  --  2.2438511 -  2.2457989
     "10111011101111011101110111011101",  --  2.2458618 -  2.2478095
     "11011101111011101110111011101110",  --  2.2478724 -  2.2498202
     "11101111011101110111011101110111",  --  2.2498830 -  2.2518308
     "01110111101110111011101110111011",  --  2.2518936 -  2.2538414
     "10111011110111011101110111011101",  --  2.2539042 -  2.2558520
     "11011101111011101110111011101110",  --  2.2559149 -  2.2578626
     "11101110111011110111011101110111",  --  2.2579255 -  2.2598733
     "01110111011101110111011110111011",  --  2.2599361 -  2.2618839
     "10111011101110111011101110111011",  --  2.2619467 -  2.2638945
     "10111101110111011101110111011101",  --  2.2639573 -  2.2659051
     "11011101110111011101111011101110",  --  2.2659679 -  2.2679157
     "11101110111011101110111011101110",  --  2.2679786 -  2.2699264
     "11101110111011101111011101110111",  --  2.2699892 -  2.2719370
     "01110111011101110111011101110111",  --  2.2719998 -  2.2739476
     "01110111011101110111011101111011",  --  2.2740104 -  2.2759582
     "10111011101110111011101110111011",  --  2.2760210 -  2.2779688
     "10111011101110111011101110111011",  --  2.2780317 -  2.2799795
     "10111011101110111011101110111011",  --  2.2800423 -  2.2819901
     "10111011101110111101110111011101",  --  2.2820529 -  2.2840007
     "11011101110111011101110111011101",  --  2.2840635 -  2.2860113
     "11011101110111011101110111011101",  --  2.2860741 -  2.2880219
     "11011101110111011101110111011101",  --  2.2880848 -  2.2900325
     "11011101110111011101110111011101",  --  2.2900954 -  2.2920432
     "11011101110111011101110111011101",  --  2.2921060 -  2.2940538
     "11011101110110111011101110111011",  --  2.2941166 -  2.2960644
     "10111011101110111011101110111011",  --  2.2961272 -  2.2980750
     "10111011101110111011101110111011",  --  2.2981379 -  2.3000856
     "10111011101110111011101110111011",  --  2.3001485 -  2.3020963
     "10110111011101110111011101110111",  --  2.3021591 -  2.3041069
     "01110111011101110111011101110111",  --  2.3041697 -  2.3061175
     "01110111011011101110111011101110",  --  2.3061803 -  2.3081281
     "11101110111011101110111011101110",  --  2.3081910 -  2.3101387
     "11101101110111011101110111011101",  --  2.3102016 -  2.3121494
     "11011101110111011101110110111011",  --  2.3122122 -  2.3141600
     "10111011101110111011101110111011",  --  2.3142228 -  2.3161706
     "10110111011101110111011101110111",  --  2.3162334 -  2.3181812
     "01110111011011101110111011101110",  --  2.3182441 -  2.3201918
     "11101110111011011101110111011101",  --  2.3202547 -  2.3222025
     "11011101110111011011101110111011",  --  2.3222653 -  2.3242131
     "10111011101110110111011101110111",  --  2.3242759 -  2.3262237
     "01110111011101101110111011101110",  --  2.3262865 -  2.3282343
     "11101110110111011101110111011101",  --  2.3282971 -  2.3302449
     "11011011101110111011101110111011",  --  2.3303078 -  2.3322556
     "01110111011101110111011101101110",  --  2.3323184 -  2.3342662
     "11101110111011101101110111011101",  --  2.3343290 -  2.3362768
     "11011101101110111011101110111011",  --  2.3363396 -  2.3382874
     "01110111011101110111011011101110",  --  2.3383502 -  2.3402980
     "11101110111011011101110111011101",  --  2.3403609 -  2.3423087
     "10111011101110111011101101110111",  --  2.3423715 -  2.3443193
     "01110111011011101110111011101101",  --  2.3443821 -  2.3463299
     "11011101110111011011101110111011",  --  2.3463927 -  2.3483405
     "10110111011101110111011011101110",  --  2.3484033 -  2.3503511
     "11101110110111011101110110111011",  --  2.3504140 -  2.3523617
     "10111011101101110111011101101110",  --  2.3524246 -  2.3543724
     "11101110111011011101110111011011",  --  2.3544352 -  2.3563830
     "10111011101110110111011101110110",  --  2.3564458 -  2.3583936
     "11101110111011011101110111011011",  --  2.3584564 -  2.3604042
     "10111011101101110111011101101110",  --  2.3604671 -  2.3624148
     "11101110110111011101110110111011",  --  2.3624777 -  2.3644255
     "10111011011101110111011011101110",  --  2.3644883 -  2.3664361
     "11101101110111011101101110111011",  --  2.3664989 -  2.3684467
     "01110111011101101110111011101101",  --  2.3685095 -  2.3704573
     "11011101101110111011101101110111",  --  2.3705202 -  2.3724679
     "01101110111011101101110111011011",  --  2.3725308 -  2.3744786
     "10111011101101110111011011101110",  --  2.3745414 -  2.3764892
     "11011101110111011011101110110111",  --  2.3765520 -  2.3784998
     "01110110111011101110110111011101",  --  2.3785626 -  2.3805104
     "10111011101101110111011011101110",  --  2.3805732 -  2.3825210
     "11011101110111011011101110110111",  --  2.3825839 -  2.3845317
     "01110110111011101101110111011011",  --  2.3845945 -  2.3865423
     "10111011011101110110111011101101",  --  2.3866051 -  2.3885529
     "11011101101110111011011101110110",  --  2.3886157 -  2.3905635
     "11101110110111011101101110111011",  --  2.3906263 -  2.3925741
     "01110110111011101101110111011011",  --  2.3926370 -  2.3945848
     "10111011011101110110111011011101",  --  2.3946476 -  2.3965954
     "11011011101110110111011101101110",  --  2.3966582 -  2.3986060
     "11011101110110111011101101110110",  --  2.3986688 -  2.4006166
     "11101110110111011101101110110111",  --  2.4006794 -  2.4026272
     "01110110111011101101110110111011",  --  2.4026901 -  2.4046378
     "10110111011011101110110111011011",  --  2.4047007 -  2.4066485
     "10111011011101101110111011011101",  --  2.4067113 -  2.4086591
     "10111011101101110110111011101101",  --  2.4087219 -  2.4106697
     "11011011101110110111011011101110",  --  2.4107325 -  2.4126803
     "11011101101110110111011101101110",  --  2.4127432 -  2.4146909
     "11011101110110111011011101101110",  --  2.4147538 -  2.4167016
     "11101101110110111011011101110110",  --  2.4167644 -  2.4187122
     "11101101110110111011011101110110",  --  2.4187750 -  2.4207228
     "11101101110110111011101101110110",  --  2.4207856 -  2.4227334
     "11101101110110111011011101110110",  --  2.4227963 -  2.4247440
     "11101101110110111011011101110110",  --  2.4248069 -  2.4267547
     "11101101110110111011011101101110",  --  2.4268175 -  2.4287653
     "11011101101110111011011101101110",  --  2.4288281 -  2.4307759
     "11011101101110110111011011101101",  --  2.4308387 -  2.4327865
     "11011011101101110111011011101101",  --  2.4328494 -  2.4347971
     "11011011101101110110111011011101",  --  2.4348600 -  2.4368078
     "10111011011101101110110111011011",  --  2.4368706 -  2.4388184
     "10110111011011101101110110111011",  --  2.4388812 -  2.4408290
     "01110110111011011101101110110111",  --  2.4408918 -  2.4428396
     "01101110110111011011101101110110",  --  2.4429024 -  2.4448502
     "11101101110110111011011101101101",  --  2.4449131 -  2.4468609
     "11011011101101110110111011011101",  --  2.4469237 -  2.4488715
     "10111011011101101110110111011011",  --  2.4489343 -  2.4508821
     "01110110111011011101101110110111",  --  2.4509449 -  2.4528927
     "01101110110110111011011101101110",  --  2.4529555 -  2.4549033
     "11011101101110110110111011011101",  --  2.4549662 -  2.4569140
     "10111011011101101101110110111011",  --  2.4569768 -  2.4589246
     "01110110111011011011101101110110",  --  2.4589874 -  2.4609352
     "11101101101110110111011011101101",  --  2.4609980 -  2.4629458
     "11011011011101101110110110111011",  --  2.4630086 -  2.4649564
     "01110110111011011011101101110110",  --  2.4650193 -  2.4669670
     "11101101101110110111011011011101",  --  2.4670299 -  2.4689777
     "10111011011011101101110110111011",  --  2.4690405 -  2.4709883
     "01101110110111011011011101101110",  --  2.4710511 -  2.4729989
     "11011011101101110110110111011011",  --  2.4730617 -  2.4750095
     "10110110111011011011101101110110",  --  2.4750724 -  2.4770201
     "11011101101110110110111011011011",  --  2.4770830 -  2.4790308
     "10110111011011011101101110110110",  --  2.4790936 -  2.4810414
     "11101101101110110110111011011101",  --  2.4811042 -  2.4830520
     "10110111011011011101101110110110",  --  2.4831148 -  2.4850626
     "11101101101110110110111011011101",  --  2.4851255 -  2.4870732
     "10110111011011011101101101110110",  --  2.4871361 -  2.4890839
     "11011101101101110110110111011011",  --  2.4891467 -  2.4910945
     "10110110111011011011101101101110",  --  2.4911573 -  2.4931051
     "11011011101101101110110110111011",  --  2.4931679 -  2.4951157
     "01101110110110111011011011101101",  --  2.4951785 -  2.4971263
     "10111011011011101101101110110110",  --  2.4971892 -  2.4991370
     "11101101101101110110110111011011",  --  2.4991998 -  2.5011476
     "01110110110111011011011101101101",  --  2.5012104 -  2.5031582
     "11011011011011101101101110110110",  --  2.5032210 -  2.5051688
     "11101101101101110110110111011011",  --  2.5052316 -  2.5071794
     "01110110110110111011011011101101",  --  2.5072423 -  2.5091901
     "10111011011011011101101101110110",  --  2.5092529 -  2.5112007
     "11011011101101101110110110110111",  --  2.5112635 -  2.5132113
     "01101101101110110110111011011011",  --  2.5132741 -  2.5152219
     "01110110110111011011011011101101",  --  2.5152847 -  2.5172325
     "10110111011011011011101101101110",  --  2.5172954 -  2.5192431
     "11011011011101101101101110110110",  --  2.5193060 -  2.5212538
     "11011101101101101110110110110111",  --  2.5213166 -  2.5232644
     "01101101101110110110110111011011",  --  2.5233272 -  2.5252750
     "01101110110110110111011011011011",  --  2.5253378 -  2.5272856
     "10110110110111011011011011011101",  --  2.5273485 -  2.5292962
     "10110110111011011011011101101101",  --  2.5293591 -  2.5313069
     "10111011011011011011101101101101",  --  2.5313697 -  2.5333175
     "11011011011011011101101101101110",  --  2.5333803 -  2.5353281
     "11011011011011101101101101101110",  --  2.5353909 -  2.5373387
     "11011011011011101101101101110110",  --  2.5374016 -  2.5393493
     "11011011011101101101101101110110",  --  2.5394122 -  2.5413600
     "11011011011101101101101101110110",  --  2.5414228 -  2.5433706
     "11011011011101101101101101101110",  --  2.5434334 -  2.5453812
     "11011011011011101101101101101110",  --  2.5454440 -  2.5473918
     "11011011011011011101101101101101",  --  2.5474547 -  2.5494024
     "11011011011011011011101101101101",  --  2.5494653 -  2.5514131
     "10110111011011011011011011101101",  --  2.5514759 -  2.5534237
     "10110110110111011011011011011011",  --  2.5534865 -  2.5554343
     "10110110110110110111011011011011",  --  2.5554971 -  2.5574449
     "01101101110110110110110110111011",  --  2.5575077 -  2.5594555
     "01101101101101101110110110110110",  --  2.5595184 -  2.5614662
     "11011011101101101101101101101110",  --  2.5615290 -  2.5634768
     "11011011011011011011101101101101",  --  2.5635396 -  2.5654874
     "10110110110111011011011011011011",  --  2.5655502 -  2.5674980
     "01110110110110110110110110111011",  --  2.5675608 -  2.5695086
     "01101101101101101101101110110110",  --  2.5695715 -  2.5715193
     "11011011011011011101101101101101",  --  2.5715821 -  2.5735299
     "10110110110111011011011011011011",  --  2.5735927 -  2.5755405
     "01101101101110110110110110110110",  --  2.5756033 -  2.5775511
     "11011011101101101101101101101101",  --  2.5776139 -  2.5795617
     "10110110111011011011011011011011",  --  2.5796246 -  2.5815723
     "01101101101110110110110110110110",  --  2.5816352 -  2.5835830
     "11011011011011101101101101101101",  --  2.5836458 -  2.5855936
     "10110110110110110110111011011011",  --  2.5856564 -  2.5876042
     "01101101101101101101101101101101",  --  2.5876670 -  2.5896148
     "11011011011011011011011011011011",  --  2.5896777 -  2.5916254
     "01101101101101101110110110110110",  --  2.5916883 -  2.5936361
     "11011011011011011011011011011011",  --  2.5936989 -  2.5956467
     "01101101110110110110110110110110",  --  2.5957095 -  2.5976573
     "11011011011011011011011011011011",  --  2.5977201 -  2.5996679
     "01101101101110110110110110110110",  --  2.5997308 -  2.6016785
     "11011011011011011011011011011011",  --  2.6017414 -  2.6036892
     "01101101101101101101101101101101",  --  2.6037520 -  2.6056998
     "10110111011011011011011011011011",  --  2.6057626 -  2.6077104
     "01101101101101101101101101101101",  --  2.6077732 -  2.6097210
     "10110110110110110110110110110110",  --  2.6097838 -  2.6117316
     "11011011011011011011011011011011",  --  2.6117945 -  2.6137423
     "01101101101101101101101101101101",  --  2.6138051 -  2.6157529
     "10110110110110110110110110110110",  --  2.6158157 -  2.6177635
     "11011011011011011011011011011011",  --  2.6178263 -  2.6197741
     "01101101101101101101101101101101",  --  2.6198369 -  2.6217847
     "10110110110110110110110110110110",  --  2.6218476 -  2.6237954
     "11011011011011011011010110110110",  --  2.6238582 -  2.6258060
     "11011011011011011011011011011011",  --  2.6258688 -  2.6278166
     "01101101101101101101101101101101",  --  2.6278794 -  2.6298272
     "10110110110110110101101101101101",  --  2.6298900 -  2.6318378
     "10110110110110110110110110110110",  --  2.6319007 -  2.6338484
     "11011011011011011011010110110110",  --  2.6339113 -  2.6358591
     "11011011011011011011011011011011",  --  2.6359219 -  2.6378697
     "01101101101011011011011011011011",  --  2.6379325 -  2.6398803
     "01101101101101101101101101011011",  --  2.6399431 -  2.6418909
     "01101101101101101101101101101101",  --  2.6419538 -  2.6439015
     "10110101101101101101101101101101",  --  2.6439644 -  2.6459122
     "10110110110101101101101101101101",  --  2.6459750 -  2.6479228
     "10110110110110101101101101101101",  --  2.6479856 -  2.6499334
     "10110110110110110101101101101101",  --  2.6499962 -  2.6519440
     "10110110110110110101101101101101",  --  2.6520069 -  2.6539546
     "10110110110110101101101101101101",  --  2.6540175 -  2.6559653
     "10110110110101101101101101101101",  --  2.6560281 -  2.6579759
     "10110101101101101101101101101101",  --  2.6580387 -  2.6599865
     "10101101101101101101101101011011",  --  2.6600493 -  2.6619971
     "01101101101101101101011011011011",  --  2.6620600 -  2.6640077
     "01101101101011011011011011011011",  --  2.6640706 -  2.6660184
     "01011011011011011011011010110110",  --  2.6660812 -  2.6680290
     "11011011011010110110110110110110",  --  2.6680918 -  2.6700396
     "11010110110110110110110101101101",  --  2.6701024 -  2.6720502
     "10110110110101101101101101101101",  --  2.6721130 -  2.6740608
     "01101101101101101101011011011011",  --  2.6741237 -  2.6760715
     "01101101011011011011011010110110",  --  2.6761343 -  2.6780821
     "11011011010110110110110110110101",  --  2.6781449 -  2.6800927
     "10110110110110101101101101101101",  --  2.6801555 -  2.6821033
     "01101101101101101011011011011011",  --  2.6821661 -  2.6841139
     "01011011011011011010110110110110",  --  2.6841768 -  2.6861246
     "11010110110110110101101101101101",  --  2.6861874 -  2.6881352
     "10101101101101101011011011011011",  --  2.6881980 -  2.6901458
     "01011011011011010110110110110110",  --  2.6902086 -  2.6921564
     "10110110110110101101101101101011",  --  2.6922192 -  2.6941670
     "01101101101011011011011010110110",  --  2.6942299 -  2.6961776
     "11011010110110110110101101101101",  --  2.6962405 -  2.6981883
     "10101101101101101011011011011010",  --  2.6982511 -  2.7001989
     "11011011011010110110110101101101",  --  2.7002617 -  2.7022095
     "10110101101101101101011011011010",  --  2.7022723 -  2.7042201
     "11011011011010110110110110101101",  --  2.7042830 -  2.7062307
     "10110101101101101101011011011010",  --  2.7062936 -  2.7082414
     "11011011010110110110110101101101",  --  2.7083042 -  2.7102520
     "10101101101101011011011011010110",  --  2.7103148 -  2.7122626
     "11011010110110110101101101101011",  --  2.7123254 -  2.7142732
     "01101101011011011010110110110110",  --  2.7143361 -  2.7162838
     "10110110110101101101101011011011",  --  2.7163467 -  2.7182945
     "01011011011010110110110101101101",  --  2.7183573 -  2.7203051
     "10101101101101011011010110110110",  --  2.7203679 -  2.7223157
     "10110110110101101101101011011011",  --  2.7223785 -  2.7243263
     "01011011011010110110101101101101",  --  2.7243891 -  2.7263369
     "01101101101011011010110110110101",  --  2.7263998 -  2.7283476
     "10110110101101101011011011010110",  --  2.7284104 -  2.7303582
     "11011010110110101101101101011011",  --  2.7304210 -  2.7323688
     "01011011011010110110101101101101",  --  2.7324316 -  2.7343794
     "01101101011011011010110110101101",  --  2.7344422 -  2.7363900
     "10110101101101011011011010110110",  --  2.7364529 -  2.7384007
     "10110110101101101101011011010110",  --  2.7384635 -  2.7404113
     "11010110110110101101101011011010",  --  2.7404741 -  2.7424219
     "11011011010110110101101101011011",  --  2.7424847 -  2.7444325
     "01011011011010110110101101101011",  --  2.7444953 -  2.7464431
     "01101011011010110110110101101101",  --  2.7465060 -  2.7484537
     "01101101011011010110110101101101",  --  2.7485166 -  2.7504644
     "01101101011011010110110101101101",  --  2.7505272 -  2.7524750
     "10101101101011011010110110101101",  --  2.7525378 -  2.7544856
     "10101101101011011010110110101101",  --  2.7545484 -  2.7564962
     "10101101101011011010110110101101",  --  2.7565591 -  2.7585068
     "10101101011011010110110101101101",  --  2.7585697 -  2.7605175
     "01101101011011010110110101101101",  --  2.7605803 -  2.7625281
     "01101101011011010110101101101011",  --  2.7625909 -  2.7645387
     "01101011011010110110101101011011",  --  2.7646015 -  2.7665493
     "01011011010110110101101101011010",  --  2.7666122 -  2.7685599
     "11011010110110101101101011010110",  --  2.7686228 -  2.7705706
     "11010110110101101101011010110110",  --  2.7706334 -  2.7725812
     "10110110101101011011010110110101",  --  2.7726440 -  2.7745918
     "10101101101011011010110101101101",  --  2.7746546 -  2.7766024
     "01101101011010110110101101101011",  --  2.7766653 -  2.7786130
     "01011011010110101101101011011010",  --  2.7786759 -  2.7806237
     "11010110110101101011011010110101",  --  2.7806865 -  2.7826343
     "10110101101101011010110110101101",  --  2.7826971 -  2.7846449
     "01101101011010110110101101011011",  --  2.7847077 -  2.7866555
     "01011010110110101101011011010110",  --  2.7867183 -  2.7886661
     "10110110101101011010110110101101",  --  2.7887290 -  2.7906768
     "01101101011010110110101101011011",  --  2.7907396 -  2.7926874
     "01011010110101101101011010110110",  --  2.7927502 -  2.7946980
     "10110101101011011010110101101101",  --  2.7947608 -  2.7967086
     "01101011010110110101101011010110",  --  2.7967714 -  2.7987192
     "11010110101101011011010110101101",  --  2.7987821 -  2.8007299
     "01101101011010110101101101011010",  --  2.8007927 -  2.8027405
     "11010110110101101011010110110101",  --  2.8028033 -  2.8047511
     "10101101011010110110101101011010",  --  2.8048139 -  2.8067617
     "11010110110101101011010110101101",  --  2.8068245 -  2.8087723
     "10101101011010110101101101011010",  --  2.8088352 -  2.8107829
     "11010110101101101011010110101101",  --  2.8108458 -  2.8127936
     "01101011011010110101101011010110",  --  2.8128564 -  2.8148042
     "10110101101101011010110101101011",  --  2.8148670 -  2.8168148
     "01011010110110101101011010110101",  --  2.8168776 -  2.8188254
     "10101101011010110110101101011010",  --  2.8188883 -  2.8208360
     "11010110101101011010110101101101",  --  2.8208989 -  2.8228467
     "01101011010110101101011010110101",  --  2.8229095 -  2.8248573
     "10101101011010110110101101011010",  --  2.8249201 -  2.8268679
     "11010110101101011010110101101011",  --  2.8269307 -  2.8288785
     "01011010110101101011010110101101",  --  2.8289414 -  2.8308891
     "01101011010110110101101011010110",  --  2.8309520 -  2.8328998
     "10110101101011010110101101011010",  --  2.8329626 -  2.8349104
     "11010110101101011010110101101011",  --  2.8349732 -  2.8369210
     "01011010110101101011010110101101",  --  2.8369838 -  2.8389316
     "01101011010101101011010110101101",  --  2.8389944 -  2.8409422
     "01101011010110101101011010110101",  --  2.8410051 -  2.8429529
     "10101101011010110101101011010110",  --  2.8430157 -  2.8449635
     "10110101011010110101101011010110",  --  2.8450263 -  2.8469741
     "10110101101011010110101101011010",  --  2.8470369 -  2.8489847
     "10110101101011010110101101011010",  --  2.8490475 -  2.8509953
     "11010110101011010110101101011010",  --  2.8510582 -  2.8530060
     "11010110101101010110101101011010",  --  2.8530688 -  2.8550166
     "11010110101101010110101101011010",  --  2.8550794 -  2.8570272
     "11010110101101010110101101011010",  --  2.8570900 -  2.8590378
     "11010110101011010110101101011010",  --  2.8591006 -  2.8610484
     "10110101101011010110101101010110",  --  2.8611113 -  2.8630590
     "10110101101011010101101011010110",  --  2.8631219 -  2.8650697
     "10110101011010110101101011010101",  --  2.8651325 -  2.8670803
     "10101101011010101101011010110101",  --  2.8671431 -  2.8690909
     "10101011010110101101010110101101",  --  2.8691537 -  2.8711015
     "01101010110101101011010101101011",  --  2.8711644 -  2.8731121
     "01011010101101011010110101011010",  --  2.8731750 -  2.8751228
     "11010110101011010110101011010110",  --  2.8751856 -  2.8771334
     "10110101011010110101011010110101",  --  2.8771962 -  2.8791440
     "10101011010110101011010110101101",  --  2.8792068 -  2.8811546
     "01011010110101011010110101011010",  --  2.8812175 -  2.8831652
     "11010110101011010110101011010110",  --  2.8832281 -  2.8851759
     "10101101011010101101011010101101",  --  2.8852387 -  2.8871865
     "01101010110101101010110101101010",  --  2.8872493 -  2.8891971
     "11010110101011010110101011010110",  --  2.8892599 -  2.8912077
     "10101101011010101101011010101101",  --  2.8912706 -  2.8932183
     "01011010110101011010110101011010",  --  2.8932812 -  2.8952290
     "11010101101010110101101010110101",  --  2.8952918 -  2.8972396
     "10101011010101101011010101101010",  --  2.8973024 -  2.8992502
     "11010110101011010101101011010101",  --  2.8993130 -  2.9012608
     "10101011010110101011010101101011",  --  2.9013236 -  2.9032714
     "01010110101011010110101011010101",  --  2.9033343 -  2.9052821
     "10101101010110101011010101101011",  --  2.9053449 -  2.9072927
     "01010110101011010101101011010101",  --  2.9073555 -  2.9093033
     "10101011010101101010110101101010",  --  2.9093661 -  2.9113139
     "11010101101010110101011010110101",  --  2.9113767 -  2.9133245
     "01101010110101011010101101010110",  --  2.9133874 -  2.9153352
     "10110101011010101101010110101011",  --  2.9153980 -  2.9173458
     "01010110101011010101101010110101",  --  2.9174086 -  2.9193564
     "10101011010101101010110101011010",  --  2.9194192 -  2.9213670
     "10110101011010101101010110101011",  --  2.9214298 -  2.9233776
     "01010110101011010101101010110101",  --  2.9234405 -  2.9253882
     "01101010110101011010101101010110",  --  2.9254511 -  2.9273989
     "10101101010110101011010101101010",  --  2.9274617 -  2.9294095
     "11010101101010101101010110101011",  --  2.9294723 -  2.9314201
     "01010110101011010101101010110101",  --  2.9314829 -  2.9334307
     "01101010110101010110101011010101",  --  2.9334936 -  2.9354413
     "10101011010101101010101101010110",  --  2.9355042 -  2.9374520
     "10101101010110101011010101011010",  --  2.9375148 -  2.9394626
     "10110101011010101101010101101010",  --  2.9395254 -  2.9414732
     "11010101101010101101010110101011",  --  2.9415360 -  2.9434838
     "01010101101010110101011010101011",  --  2.9435467 -  2.9454944
     "01010110101011010101011010101101",  --  2.9455573 -  2.9475051
     "01010110101011010101101010101101",  --  2.9475679 -  2.9495157
     "01011010101011010101101010101101",  --  2.9495785 -  2.9515263
     "01011010101011010101101010101101",  --  2.9515891 -  2.9535369
     "01011010101011010101101010101101",  --  2.9535997 -  2.9555475
     "01011010101011010101011010101101",  --  2.9556104 -  2.9575582
     "01010110101011010101011010101011",  --  2.9576210 -  2.9595688
     "01010110101010110101010110101011",  --  2.9596316 -  2.9615794
     "01010101101010101101010101101010",  --  2.9616422 -  2.9635900
     "11010101011010101011010101011010",  --  2.9636528 -  2.9656006
     "10101101010110101010110101010110",  --  2.9656635 -  2.9676113
     "10101011010101011010101011010101",  --  2.9676741 -  2.9696219
     "10101010110101010110101010110101",  --  2.9696847 -  2.9716325
     "01011010101011010101011010101011",  --  2.9716953 -  2.9736431
     "01010101101010101101010101101010",  --  2.9737059 -  2.9756537
     "10110101010110101010110101010101",  --  2.9757166 -  2.9776643
     "10101010110101010110101010110101",  --  2.9777272 -  2.9796750
     "01011010101011010101010110101010",  --  2.9797378 -  2.9816856
     "11010101011010101011010101010110",  --  2.9817484 -  2.9836962
     "10101011010101011010101011010101",  --  2.9837590 -  2.9857068
     "01011010101011010101010110101010",  --  2.9857697 -  2.9877174
     "11010101011010101010110101010110",  --  2.9877803 -  2.9897281
     "10101010110101010110101010101101",  --  2.9897909 -  2.9917387
     "01010110101010101101010101011010",  --  2.9918015 -  2.9937493
     "10101101010101011010101011010101",  --  2.9938121 -  2.9957599
     "01011010101010110101010101101010",  --  2.9958228 -  2.9977705
     "10110101010101101010101011010101",  --  2.9978334 -  2.9997812
     "01011010101010110101010110101010",  --  2.9998440 -  3.0017918
     "10110101010101101010101011010101",  --  3.0018546 -  3.0038024
     "01011010101010110101010101101010",  --  3.0038652 -  3.0058130
     "10101101010101011010101010110101",  --  3.0058759 -  3.0078236
     "01010101101010101011010101010110",  --  3.0078865 -  3.0098343
     "10101010110101010101011010101010",  --  3.0098971 -  3.0118449
     "11010101010110101010101011010101",  --  3.0119077 -  3.0138555
     "01011010101010110101010101011010",  --  3.0139183 -  3.0158661
     "10101011010101010101101010101011",  --  3.0159289 -  3.0178767
     "01010101010110101010101011010101",  --  3.0179396 -  3.0198874
     "01011010101010101101010101010110",  --  3.0199502 -  3.0218980
     "10101010101101010101010110101010",  --  3.0219608 -  3.0239086
     "10101101010101010110101010101011",  --  3.0239714 -  3.0259192
     "01010101010110101010101011010101",  --  3.0259820 -  3.0279298
     "01010110101010101011010101010101",  --  3.0279927 -  3.0299405
     "10101010101010110101010101011010",  --  3.0300033 -  3.0319511
     "10101010110101010101010110101010",  --  3.0320139 -  3.0339617
     "10101101010101010101101010101010",  --  3.0340245 -  3.0359723
     "11010101010101011010101010101011",  --  3.0360351 -  3.0379829
     "01010101010101101010101010110101",  --  3.0380458 -  3.0399935
     "01010101011010101010101011010101",  --  3.0400564 -  3.0420042
     "01010101011010101010101011010101",  --  3.0420670 -  3.0440148
     "01010101101010101010101101010101",  --  3.0440776 -  3.0460254
     "01010101101010101010101101010101",  --  3.0460882 -  3.0480360
     "01010101101010101010101101010101",  --  3.0480989 -  3.0500466
     "01010101101010101010101011010101",  --  3.0501095 -  3.0520573
     "01010101011010101010101010110101",  --  3.0521201 -  3.0540679
     "01010101010110101010101010101101",  --  3.0541307 -  3.0560785
     "01010101010101011010101010101010",  --  3.0561413 -  3.0580891
     "11010101010101010101101010101010",  --  3.0581520 -  3.0600997
     "10101101010101010101010110101010",  --  3.0601626 -  3.0621104
     "10101010101101010101010101010110",  --  3.0621732 -  3.0641210
     "10101010101010101011010101010101",  --  3.0641838 -  3.0661316
     "01010110101010101010101010110101",  --  3.0661944 -  3.0681422
     "01010101010101011010101010101010",  --  3.0682050 -  3.0701528
     "10110101010101010101010101101010",  --  3.0702157 -  3.0721635
     "10101010101010110101010101010101",  --  3.0722263 -  3.0741741
     "01010110101010101010101010101101",  --  3.0742369 -  3.0761847
     "01010101010101010101101010101010",  --  3.0762475 -  3.0781953
     "10101010101101010101010101010101",  --  3.0782581 -  3.0802059
     "01011010101010101010101010101101",  --  3.0802688 -  3.0822166
     "01010101010101010101011010101010",  --  3.0822794 -  3.0842272
     "10101010101010101101010101010101",  --  3.0842900 -  3.0862378
     "01010101010110101010101010101010",  --  3.0863006 -  3.0882484
     "10101011010101010101010101010101",  --  3.0883112 -  3.0902590
     "01011010101010101010101010101010",  --  3.0903219 -  3.0922696
     "10110101010101010101010101010101",  --  3.0923325 -  3.0942803
     "01101010101010101010101010101010",  --  3.0943431 -  3.0962909
     "10110101010101010101010101010101",  --  3.0963537 -  3.0983015
     "01011010101010101010101010101010",  --  3.0983643 -  3.1003121
     "10101010110101010101010101010101",  --  3.1003750 -  3.1023227
     "01010101010101101010101010101010",  --  3.1023856 -  3.1043334
     "10101010101010101010101101010101",  --  3.1043962 -  3.1063440
     "01010101010101010101010101010101",  --  3.1064068 -  3.1083546
     "01101010101010101010101010101010",  --  3.1084174 -  3.1103652
     "10101010101010101011010101010101",  --  3.1104281 -  3.1123758
     "01010101010101010101010101010101",  --  3.1124387 -  3.1143865
     "01010101101010101010101010101010",  --  3.1144493 -  3.1163971
     "10101010101010101010101010101010",  --  3.1164599 -  3.1184077
     "10101101010101010101010101010101",  --  3.1184705 -  3.1204183
     "01010101010101010101010101010101",  --  3.1204812 -  3.1224289
     "01010101010101101010101010101010",  --  3.1224918 -  3.1244396
     "10101010101010101010101010101010",  --  3.1245024 -  3.1264502
     "10101010101010101010101010101010",  --  3.1265130 -  3.1284608
     "10101010101010101101010101010101",  --  3.1285236 -  3.1304714
     "01010101010101010101010101010101",  --  3.1305342 -  3.1324820
     "01010101010101010101010101010101",  --  3.1325449 -  3.1344927
     "01010101010101010101010101010101",  --  3.1345555 -  3.1365033
     "01010101010101010101010101010101",  --  3.1365661 -  3.1385139
     "01010101010101010101010101010101",  --  3.1385767 -  3.1405245
     "01010101010101010101010101010101",  --  3.1405873 -  3.1425351
     "01010101010101010101010101010101",  --  3.1425980 -  3.1445458
     "01010101010101010101010101010101",  --  3.1446086 -  3.1465564
     "01010101010101010101010101010101",  --  3.1466192 -  3.1485670
     "01010101010101010101010101010101",  --  3.1486298 -  3.1505776
     "01010101010101010101010101010101",  --  3.1506404 -  3.1525882
     "01010101010101010010101010101010",  --  3.1526511 -  3.1545988
     "10101010101010101010101010101010",  --  3.1546617 -  3.1566095
     "10101010101010101010101010101010",  --  3.1566723 -  3.1586201
     "10101010101010101010010101010101",  --  3.1586829 -  3.1606307
     "01010101010101010101010101010101",  --  3.1606935 -  3.1626413
     "01010101010101010101010101010010",  --  3.1627042 -  3.1646519
     "10101010101010101010101010101010",  --  3.1647148 -  3.1666626
     "10101010101010101010101010010101",  --  3.1667254 -  3.1686732
     "01010101010101010101010101010101",  --  3.1687360 -  3.1706838
     "01010101010101001010101010101010",  --  3.1707466 -  3.1726944
     "10101010101010101010101010101010",  --  3.1727573 -  3.1747050
     "01010101010101010101010101010101",  --  3.1747679 -  3.1767157
     "01010101010010101010101010101010",  --  3.1767785 -  3.1787263
     "10101010101010101010010101010101",  --  3.1787891 -  3.1807369
     "01010101010101010101010100101010",  --  3.1807997 -  3.1827475
     "10101010101010101010101010101001",  --  3.1828103 -  3.1847581
     "01010101010101010101010101010100",  --  3.1848210 -  3.1867688
     "10101010101010101010101010101010",  --  3.1868316 -  3.1887794
     "01010101010101010101010101010100",  --  3.1888422 -  3.1907900
     "10101010101010101010101010101001",  --  3.1908528 -  3.1928006
     "01010101010101010101010101001010",  --  3.1928634 -  3.1948112
     "10101010101010101010100101010101",  --  3.1948741 -  3.1968219
     "01010101010101010010101010101010",  --  3.1968847 -  3.1988325
     "10101010101001010101010101010101",  --  3.1988953 -  3.2008431
     "01010010101010101010101010101001",  --  3.2009059 -  3.2028537
     "01010101010101010101010010101010",  --  3.2029165 -  3.2048643
     "10101010101010010101010101010101",  --  3.2049272 -  3.2068749
     "01010010101010101010101010100101",  --  3.2069378 -  3.2088856
     "01010101010101010100101010101010",  --  3.2089484 -  3.2108962
     "10101010010101010101010101010100",  --  3.2109590 -  3.2129068
     "10101010101010101001010101010101",  --  3.2129696 -  3.2149174
     "01010100101010101010101010100101",  --  3.2149803 -  3.2169280
     "01010101010101001010101010101010",  --  3.2169909 -  3.2189387
     "10100101010101010101010010101010",  --  3.2190015 -  3.2209493
     "10101010100101010101010101010010",  --  3.2210121 -  3.2229599
     "10101010101010010101010101010101",  --  3.2230227 -  3.2249705
     "00101010101010101001010101010101",  --  3.2250334 -  3.2269811
     "01010010101010101010100101010101",  --  3.2270440 -  3.2289918
     "01010100101010101010101001010101",  --  3.2290546 -  3.2310024
     "01010101001010101010101010010101",  --  3.2310652 -  3.2330130
     "01010101010010101010101010010101",  --  3.2330758 -  3.2350236
     "01010101010010101010101010010101",  --  3.2350865 -  3.2370342
     "01010101010010101010101010010101",  --  3.2370971 -  3.2390449
     "01010101001010101010101001010101",  --  3.2391077 -  3.2410555
     "01010101001010101010101001010101",  --  3.2411183 -  3.2430661
     "01010100101010101010010101010101",  --  3.2431289 -  3.2450767
     "01001010101010101001010101010101",  --  3.2451395 -  3.2470873
     "00101010101010010101010101010010",  --  3.2471502 -  3.2490980
     "10101010100101010101010100101010",  --  3.2491608 -  3.2511086
     "10101001010101010100101010101010",  --  3.2511714 -  3.2531192
     "10010101010101001010101010100101",  --  3.2531820 -  3.2551298
     "01010101001010101010100101010101",  --  3.2551926 -  3.2571404
     "01001010101010100101010101010010",  --  3.2572033 -  3.2591511
     "10101010100101010101010010101010",  --  3.2592139 -  3.2611617
     "10100101010101010010101010101001",  --  3.2612245 -  3.2631723
     "01010101001010101010100101010101",  --  3.2632351 -  3.2651829
     "01001010101010010101010101001010",  --  3.2652457 -  3.2671935
     "10101001010101010100101010101001",  --  3.2672564 -  3.2692041
     "01010101001010101010100101010101",  --  3.2692670 -  3.2712148
     "00101010101001010101010100101010",  --  3.2712776 -  3.2732254
     "10100101010101001010101010010101",  --  3.2732882 -  3.2752360
     "01010100101010101001010101010010",  --  3.2752988 -  3.2772466
     "10101010010101010100101010101001",  --  3.2773095 -  3.2792572
     "01010101001010101010010101010100",  --  3.2793201 -  3.2812679
     "10101010100101010100101010101001",  --  3.2813307 -  3.2832785
     "01010101001010101010010101010100",  --  3.2833413 -  3.2852891
     "10101010010101010100101010101001",  --  3.2853519 -  3.2872997
     "01010101001010101001010101010010",  --  3.2873626 -  3.2893103
     "10101001010101010010101010100101",  --  3.2893732 -  3.2913210
     "01010010101010100101010100101010",  --  3.2913838 -  3.2933316
     "10100101010100101010101001010101",  --  3.2933944 -  3.2953422
     "00101010100101010101001010101001",  --  3.2954050 -  3.2973528
     "01010101001010101001010101001010",  --  3.2974156 -  3.2993634
     "10100101010101001010101001010101",  --  3.2994263 -  3.3013741
     "00101010100101010101001010101001",  --  3.3014369 -  3.3033847
     "01010100101010100101010100101010",  --  3.3034475 -  3.3053953
     "10010101010100101010100101010100",  --  3.3054581 -  3.3074059
     "10101010010101010010101010010101",  --  3.3074687 -  3.3094165
     "01001010101001010101001010101001",  --  3.3094794 -  3.3114272
     "01010100101010100101010100101010",  --  3.3114900 -  3.3134378
     "10010101001010101001010101001010",  --  3.3135006 -  3.3154484
     "10100101010100101010100101010010",  --  3.3155112 -  3.3174590
     "10101001010101001010101001010101",  --  3.3175218 -  3.3194696
     "00101010010101010010101010010101",  --  3.3195325 -  3.3214802
     "01001010100101010100101010100101",  --  3.3215431 -  3.3234909
     "01001010101001010101001010100101",  --  3.3235537 -  3.3255015
     "01010010101001010101001010101001",  --  3.3255643 -  3.3275121
     "01010010101010010101001010101001",  --  3.3275749 -  3.3295227
     "01010010101010010101001010101001",  --  3.3295856 -  3.3315333
     "01010010101010010101001010101001",  --  3.3315962 -  3.3335440
     "01010010101010010101001010100101",  --  3.3336068 -  3.3355546
     "01010010101001010101001010100101",  --  3.3356174 -  3.3375652
     "01001010101001010100101010010101",  --  3.3376280 -  3.3395758
     "01001010100101010010101010010101",  --  3.3396387 -  3.3415864
     "00101010010101010010101001010100",  --  3.3416493 -  3.3435971
     "10101001010101001010100101010010",  --  3.3436599 -  3.3456077
     "10100101010010101010010101001010",  --  3.3456705 -  3.3476183
     "10010101001010100101010100101010",  --  3.3476811 -  3.3496289
     "01010100101010010101001010100101",  --  3.3496918 -  3.3516395
     "01001010100101010010101010010101",  --  3.3517024 -  3.3536502
     "00101010010101001010100101010010",  --  3.3537130 -  3.3556608
     "10100101010010101001010100101010",  --  3.3557236 -  3.3576714
     "01010100101010010101001010100101",  --  3.3577342 -  3.3596820
     "01001010100101010010101001010100",  --  3.3597448 -  3.3616926
     "10101001010100101010010101001010",  --  3.3617555 -  3.3637033
     "10010100101010010101001010100101",  --  3.3637661 -  3.3657139
     "01001010100101010010101001010100",  --  3.3657767 -  3.3677245
     "10100101010010101001010100101010",  --  3.3677873 -  3.3697351
     "01010100101001010100101010010101",  --  3.3697979 -  3.3717457
     "00101010010100101010010101001010",  --  3.3718086 -  3.3737564
     "10010101001010010101001010100101",  --  3.3738192 -  3.3757670
     "01001010010101001010100101010010",  --  3.3758298 -  3.3777776
     "10010101001010100101001010100101",  --  3.3778404 -  3.3797882
     "01001010010101001010100101001010",  --  3.3798510 -  3.3817988
     "10010101001010010101001010100101",  --  3.3818617 -  3.3838094
     "00101010010101001010010101001010",  --  3.3838723 -  3.3858201
     "10010100101010010100101010010101",  --  3.3858829 -  3.3878307
     "00101001010100101001010100101001",  --  3.3878935 -  3.3898413
     "01010010101001010010101001010010",  --  3.3899041 -  3.3918519
     "10100101001010100101001010100101",  --  3.3919148 -  3.3938625
     "00101010010100101010010100101010",  --  3.3939254 -  3.3958732
     "01010010101001010010101001010010",  --  3.3959360 -  3.3978838
     "10100101001010100101001010100101",  --  3.3979466 -  3.3998944
     "00101001010100101001010100101001",  --  3.3999572 -  3.4019050
     "01010010100101001010100101001010",  --  3.4019679 -  3.4039156
     "10010100101001010100101001010100",  --  3.4039785 -  3.4059263
     "10100101001010100101001010100101",  --  3.4059891 -  3.4079369
     "00101001010100101001010010101001",  --  3.4079997 -  3.4099475
     "01001010010101001010010100101010",  --  3.4100103 -  3.4119581
     "01010010100101010010100101001010",  --  3.4120209 -  3.4139687
     "10010100101001010010101001010010",  --  3.4140316 -  3.4159794
     "10010101001010010100101001010100",  --  3.4160422 -  3.4179900
     "10100101001010010101001010010100",  --  3.4180528 -  3.4200006
     "10100101010010100101001010010100",  --  3.4200634 -  3.4220112
     "10101001010010100101001010100101",  --  3.4220740 -  3.4240218
     "00101001010010100101010010100101",  --  3.4240847 -  3.4260325
     "00101001010010100101010010100101",  --  3.4260953 -  3.4280431
     "00101001010010100101010010100101",  --  3.4281059 -  3.4300537
     "00101001010010100101001010100101",  --  3.4301165 -  3.4320643
     "00101001010010100101001010010100",  --  3.4321271 -  3.4340749
     "10101001010010100101001010010100",  --  3.4341378 -  3.4360855
     "10100101001010010100101001010100",  --  3.4361484 -  3.4380962
     "10100101001010010100101001010010",  --  3.4381590 -  3.4401068
     "10010100101001010010100101001010",  --  3.4401696 -  3.4421174
     "01010010100101001010010101001010",  --  3.4421802 -  3.4441280
     "01010010100101001010010100101001",  --  3.4441909 -  3.4461386
     "01001010010100101001010010100101",  --  3.4462015 -  3.4481493
     "00101001010010100101001010010100",  --  3.4482121 -  3.4501599
     "10100101001010010100100101001010",  --  3.4502227 -  3.4521705
     "01010010100101001010010100101001",  --  3.4522333 -  3.4541811
     "01001010010100101001010010100101",  --  3.4542440 -  3.4561917
     "00101001010010100100101001010010",  --  3.4562546 -  3.4582024
     "10010100101001010010100101001010",  --  3.4582652 -  3.4602130
     "01010010010100101001010010100101",  --  3.4602758 -  3.4622236
     "00101001010010100100101001010010",  --  3.4622864 -  3.4642342
     "10010100101001010010100100101001",  --  3.4642971 -  3.4662448
     "01001010010100101001010010010100",  --  3.4663077 -  3.4682555
     "10100101001010010100101001001010",  --  3.4683183 -  3.4702661
     "01010010100101001010010010100101",  --  3.4703289 -  3.4722767
     "00101001010010010100101001010010",  --  3.4723395 -  3.4742873
     "10010010100101001010010100100101",  --  3.4743501 -  3.4762979
     "00101001010010100100101001010010",  --  3.4763608 -  3.4783086
     "10010100100101001010010100100101",  --  3.4783714 -  3.4803192
     "00101001010010010100101001010010",  --  3.4803820 -  3.4823298
     "01010010100101001001010010100101",  --  3.4823926 -  3.4843404
     "00100101001010010100100101001010",  --  3.4844032 -  3.4863510
     "01010010010100101001001010010100",  --  3.4864139 -  3.4883617
     "10100100101001010010010100101001",  --  3.4884245 -  3.4903723
     "01001001010010100100101001010010",  --  3.4904351 -  3.4923829
     "01010010100100101001010010100100",  --  3.4924457 -  3.4943935
     "10100101001001010010100100101001",  --  3.4944563 -  3.4964041
     "01001001010010100100101001010010",  --  3.4964670 -  3.4984147
     "01010010100100101001010010010100",  --  3.4984776 -  3.5004254
     "10010100101001001010010100100101",  --  3.5004882 -  3.5024360
     "00101001001010010010100101001001",  --  3.5024988 -  3.5044466
     "01001010010010100100101001010010",  --  3.5045094 -  3.5064572
     "01010010010100101001001010010010",  --  3.5065201 -  3.5084678
     "10010100100101001001010010100100",  --  3.5085307 -  3.5104785
     "10100100101001010010010100100101",  --  3.5105413 -  3.5124891
     "00100101001010010010100100101001",  --  3.5125519 -  3.5144997
     "00101001010010010100100101001001",  --  3.5145625 -  3.5165103
     "01001001010010100100101001001010",  --  3.5165732 -  3.5185209
     "01001010010010100101001001010010",  --  3.5185838 -  3.5205316
     "01010010010100100101001001010010",  --  3.5205944 -  3.5225422
     "01010010010100100101001001010010",  --  3.5226050 -  3.5245528
     "10010010100100101001001010010010",  --  3.5246156 -  3.5265634
     "10010010100100101001001010010010",  --  3.5266262 -  3.5285740
     "10010010100100101001001010010010",  --  3.5286369 -  3.5305847
     "10010010010100100101001001010010",  --  3.5306475 -  3.5325953
     "01010010010100100101001001010010",  --  3.5326581 -  3.5346059
     "01010010010100100100101001001010",  --  3.5346687 -  3.5366165
     "01001010010010100100101001001001",  --  3.5366793 -  3.5386271
     "01001001010010010100100101001001",  --  3.5386900 -  3.5406378
     "00101001001010010010100100100101",  --  3.5407006 -  3.5426484
     "00100101001001010010010010100100",  --  3.5427112 -  3.5446590
     "10100100101001001001010010010100",  --  3.5447218 -  3.5466696
     "10010010100100101001001001010010",  --  3.5467324 -  3.5486802
     "01010010010010100100101001001001",  --  3.5487431 -  3.5506908
     "01001001010010010010100100101001",  --  3.5507537 -  3.5527015
     "00100101001001001010010010100100",  --  3.5527643 -  3.5547121
     "10010100100100101001001010010010",  --  3.5547749 -  3.5567227
     "01010010010010100100101001001001",  --  3.5567855 -  3.5587333
     "01001001001010010010010100100100",  --  3.5587962 -  3.5607439
     "10100100100101001001010010010010",  --  3.5608068 -  3.5627546
     "10010010010100100100101001001001",  --  3.5628174 -  3.5647652
     "01001001001010010010010100100100",  --  3.5648280 -  3.5667758
     "10100100100100101001001001010010",  --  3.5668386 -  3.5687864
     "01001010010010010100100100101001",  --  3.5688493 -  3.5707970
     "00100101001001001001010010010010",  --  3.5708599 -  3.5728077
     "10010010010100100100100101001001",  --  3.5728705 -  3.5748183
     "00101001001001010010010010010100",  --  3.5748811 -  3.5768289
     "10010010100100100100101001001001",  --  3.5768917 -  3.5788395
     "00101001001001010010010010010100",  --  3.5789024 -  3.5808501
     "10010010010100100100101001001001",  --  3.5809130 -  3.5828608
     "00101001001001001010010010010010",  --  3.5829236 -  3.5848714
     "10010010010010100100100100101001",  --  3.5849342 -  3.5868820
     "00100100101001001001001010010010",  --  3.5869448 -  3.5888926
     "01001010010010010010100100100100",  --  3.5889554 -  3.5909032
     "10100100100100100101001001001001",  --  3.5909661 -  3.5929139
     "01001001001001001010010010010010",  --  3.5929767 -  3.5949245
     "10010010010010010100100100100101",  --  3.5949873 -  3.5969351
     "00100100100100101001001001001001",  --  3.5969979 -  3.5989457
     "01001001001001001010010010010010",  --  3.5990085 -  3.6009563
     "01010010010010010010100100100100",  --  3.6010192 -  3.6029670
     "10010100100100100100100101001001",  --  3.6030298 -  3.6049776
     "00100100101001001001001001010010",  --  3.6050404 -  3.6069882
     "01001001001001010010010010010010",  --  3.6070510 -  3.6089988
     "01010010010010010010010100100100",  --  3.6090616 -  3.6110094
     "10010010010100100100100100100101",  --  3.6110723 -  3.6130200
     "00100100100100100100101001001001",  --  3.6130829 -  3.6150307
     "00100100101001001001001001001001",  --  3.6150935 -  3.6170413
     "01001001001001001001001010010010",  --  3.6171041 -  3.6190519
     "01001001001001010010010010010010",  --  3.6191147 -  3.6210625
     "01001001010010010010010010010010",  --  3.6211254 -  3.6230731
     "10010010010010010010010010010100",  --  3.6231360 -  3.6250838
     "10010010010010010010010100100100",  --  3.6251466 -  3.6270944
     "10010010010010010010100100100100",  --  3.6271572 -  3.6291050
     "10010010010010010100100100100100",  --  3.6291678 -  3.6311156
     "10010010010010010100100100100100",  --  3.6311785 -  3.6331262
     "10010010010010010010100100100100",  --  3.6331891 -  3.6351369
     "10010010010010010010010100100100",  --  3.6351997 -  3.6371475
     "10010010010010010010010010010100",  --  3.6372103 -  3.6391581
     "10010010010010010010010010010010",  --  3.6392209 -  3.6411687
     "01001001010010010010010010010010",  --  3.6412315 -  3.6431793
     "01001001001001001001001010010010",  --  3.6432422 -  3.6451900
     "01001001001001001001001001001001",  --  3.6452528 -  3.6472006
     "00100100100101001001001001001001",  --  3.6472634 -  3.6492112
     "00100100100100100100100100100100",  --  3.6492740 -  3.6512218
     "10010010010010010100100100100100",  --  3.6512846 -  3.6532324
     "10010010010010010010010010010010",  --  3.6532953 -  3.6552431
     "01001001001001001001001001001001",  --  3.6553059 -  3.6572537
     "00100100100101001001001001001001",  --  3.6573165 -  3.6592643
     "00100100100100100100100100100100",  --  3.6593271 -  3.6612749
     "10010010010010010010010010010010",  --  3.6613377 -  3.6632855
     "01001001001001001001001001001001",  --  3.6633484 -  3.6652961
     "00100100100100100100100100100100",  --  3.6653590 -  3.6673068
     "10010010010010010010010010010010",  --  3.6673696 -  3.6693174
     "01001001001001001001001001001001",  --  3.6693802 -  3.6713280
     "00100100100100100100100100100100",  --  3.6713908 -  3.6733386
     "10010010010010010010010010010010",  --  3.6734015 -  3.6753492
     "01001001001001001001001001000100",  --  3.6754121 -  3.6773599
     "10010010010010010010010010010010",  --  3.6774227 -  3.6793705
     "01001001001001001001001001001001",  --  3.6794333 -  3.6813811
     "00100100100100100100100010010010",  --  3.6814439 -  3.6833917
     "01001001001001001001001001001001",  --  3.6834546 -  3.6854023
     "00100100100100100100100100010010",  --  3.6854652 -  3.6874130
     "01001001001001001001001001001001",  --  3.6874758 -  3.6894236
     "00100100100100100010010010010010",  --  3.6894864 -  3.6914342
     "01001001001001001001001001001001",  --  3.6914970 -  3.6934448
     "00010010010010010010010010010010",  --  3.6935077 -  3.6954554
     "01001001001000100100100100100100",  --  3.6955183 -  3.6974661
     "10010010010010010010001001001001",  --  3.6975289 -  3.6994767
     "00100100100100100100100010010010",  --  3.6995395 -  3.7014873
     "01001001001001001001001000100100",  --  3.7015501 -  3.7034979
     "10010010010010010010010010001001",  --  3.7035607 -  3.7055085
     "00100100100100100100100100010010",  --  3.7055714 -  3.7075192
     "01001001001001001001000100100100",  --  3.7075820 -  3.7095298
     "10010010010010010001001001001001",  --  3.7095926 -  3.7115404
     "00100100100010010010010010010010",  --  3.7116032 -  3.7135510
     "01001000100100100100100100100100",  --  3.7136138 -  3.7155616
     "01001001001001001001000100100100",  --  3.7156245 -  3.7175723
     "10010010010010001001001001001001",  --  3.7176351 -  3.7195829
     "00100010010010010010010010001001",  --  3.7196457 -  3.7215935
     "00100100100100100010010010010010",  --  3.7216563 -  3.7236041
     "01001000100100100100100100010010",  --  3.7236669 -  3.7256147
     "01001001001001000100100100100100",  --  3.7256776 -  3.7276253
     "10001001001001001001000100100100",  --  3.7276882 -  3.7296360
     "10010010001001001001001001000100",  --  3.7296988 -  3.7316466
     "10010010010010001001001001001001",  --  3.7317094 -  3.7336572
     "00010010010010010001001001001001",  --  3.7337200 -  3.7356678
     "00100010010010010010001001001001",  --  3.7357307 -  3.7376784
     "00100010010010010010010001001001",  --  3.7377413 -  3.7396891
     "00100100010010010010010001001001",  --  3.7397519 -  3.7416997
     "00100100010010010010010001001001",  --  3.7417625 -  3.7437103
     "00100100010010010010001001001001",  --  3.7437731 -  3.7457209
     "00100010010010010010001001001001",  --  3.7457838 -  3.7477315
     "00100010010010010001001001001001",  --  3.7477944 -  3.7497422
     "00010010010010001001001001001000",  --  3.7498050 -  3.7517528
     "10010010010001001001001000100100",  --  3.7518156 -  3.7537634
     "10010001001001001001000100100100",  --  3.7538262 -  3.7557740
     "10001001001001000100100100100010",  --  3.7558368 -  3.7577846
     "01001001000100100100100010010010",  --  3.7578475 -  3.7597953
     "01000100100100100010010010010001",  --  3.7598581 -  3.7618059
     "00100100100010010010010001001001",  --  3.7618687 -  3.7638165
     "00100010010010001001001001000100",  --  3.7638793 -  3.7658271
     "10010010001001001001000100100100",  --  3.7658899 -  3.7678377
     "01001001001000100100100010010010",  --  3.7679006 -  3.7698484
     "01000100100100100010010010001001",  --  3.7699112 -  3.7718590
     "00100100010010010001001001001000",  --  3.7719218 -  3.7738696
     "10010010001001001000100100100100",  --  3.7739324 -  3.7758802
     "01001001000100100100010010010010",  --  3.7759430 -  3.7778908
     "00100100100010010010001001001001",  --  3.7779537 -  3.7799014
     "00010010010001001001000100100100",  --  3.7799643 -  3.7819121
     "01001001000100100100010010010010",  --  3.7819749 -  3.7839227
     "00100100100010010010001001001000",  --  3.7839855 -  3.7859333
     "10010010001001001000100100100010",  --  3.7859961 -  3.7879439
     "01001000100100100010010010001001",  --  3.7880068 -  3.7899545
     "00100010010010001001001000100100",  --  3.7900174 -  3.7919652
     "10001001000100100100010010010001",  --  3.7920280 -  3.7939758
     "00100100010010010001001001000100",  --  3.7940386 -  3.7959864
     "10010001001000100100100010010010",  --  3.7960492 -  3.7979970
     "00100100100010010001001001000100",  --  3.7980599 -  3.8000076
     "10010001001000100100100010010010",  --  3.8000705 -  3.8020183
     "00100100100010010001001001000100",  --  3.8020811 -  3.8040289
     "10001001001000100100100010010001",  --  3.8040917 -  3.8060395
     "00100100010010001001001000100100",  --  3.8061023 -  3.8080501
     "10001001000100100100010010001001",  --  3.8081130 -  3.8100607
     "00100010010001001001000100100010",  --  3.8101236 -  3.8120714
     "01001000100100010010001001001000",  --  3.8121342 -  3.8140820
     "10010001001001000100100010010010",  --  3.8141448 -  3.8160926
     "00100100010010001001001000100100",  --  3.8161554 -  3.8181032
     "01001000100100100010010001001001",  --  3.8181660 -  3.8201138
     "00010010001001000100100010010010",  --  3.8201767 -  3.8221245
     "00100100010010001001001000100100",  --  3.8221873 -  3.8241351
     "01001000100100010010010001001000",  --  3.8241979 -  3.8261457
     "10010001001000100100100010010001",  --  3.8262085 -  3.8281563
     "00100010010001001000100100100010",  --  3.8282191 -  3.8301669
     "01000100100010010001001000100100",  --  3.8302298 -  3.8321776
     "01001001000100100010010001001000",  --  3.8322404 -  3.8341882
     "10010001001000100100010010001001",  --  3.8342510 -  3.8361988
     "00010010010001001000100100010010",  --  3.8362616 -  3.8382094
     "00100100010010001001000100100010",  --  3.8382722 -  3.8402200
     "01000100100010010001001000100100",  --  3.8402829 -  3.8422306
     "01001000100100010010001001000100",  --  3.8422935 -  3.8442413
     "10001001000100100010010001001000",  --  3.8443041 -  3.8462519
     "10010001001000100100010010001001",  --  3.8463147 -  3.8482625
     "00010010001001000100010010001001",  --  3.8483253 -  3.8502731
     "00010010001001000100100010010001",  --  3.8503360 -  3.8522837
     "00100010010001001000100010010001",  --  3.8523466 -  3.8542944
     "00100010010001001000100100010010",  --  3.8543572 -  3.8563050
     "00100100010001001000100100010010",  --  3.8563678 -  3.8583156
     "00100100010001001000100100010010",  --  3.8583784 -  3.8603262
     "00100100010010001000100100010010",  --  3.8603891 -  3.8623368
     "00100100010001001000100100010010",  --  3.8623997 -  3.8643475
     "00100100010001001000100100010010",  --  3.8644103 -  3.8663581
     "00100010010001001000100100010001",  --  3.8664209 -  3.8683687
     "00100010010001000100100010010001",  --  3.8684315 -  3.8703793
     "00100010001001000100100010001001",  --  3.8704421 -  3.8723899
     "00010010001000100100010010001000",  --  3.8724528 -  3.8744006
     "10010001001000100010010001001000",  --  3.8744634 -  3.8764112
     "10001001000100100010001001000100",  --  3.8764740 -  3.8784218
     "10001000100100010010001000100100",  --  3.8784846 -  3.8804324
     "01000100100010010001000100100010",  --  3.8804952 -  3.8824430
     "00100100010010001000100100010001",  --  3.8825059 -  3.8844537
     "00100010010001000100100010001001",  --  3.8845165 -  3.8864643
     "00010001001000100100010001001000",  --  3.8865271 -  3.8884749
     "10001001000100010010001000100100",  --  3.8885377 -  3.8904855
     "01001000100010010001000100100010",  --  3.8905483 -  3.8924961
     "00100100010001001000100010010001",  --  3.8925590 -  3.8945067
     "00010010001000100100010001001000",  --  3.8945696 -  3.8965174
     "10001001000100010010001000100100",  --  3.8965802 -  3.8985280
     "01000100100010001001000100010001",  --  3.8985908 -  3.9005386
     "00100010001001000100010010001000",  --  3.9006014 -  3.9025492
     "10010001000100100010001000100100",  --  3.9026121 -  3.9045598
     "01000100100010001001000100010001",  --  3.9046227 -  3.9065705
     "00100010001001000100010010001000",  --  3.9066333 -  3.9085811
     "10001001000100010010001000100010",  --  3.9086439 -  3.9105917
     "01000100010010001000100010010001",  --  3.9106545 -  3.9126023
     "00010010001000100010010001000100",  --  3.9126652 -  3.9146129
     "01001000100010010001000100010010",  --  3.9146758 -  3.9166236
     "00100010001001000100010001001000",  --  3.9166864 -  3.9186342
     "10001000100100010001000100100010",  --  3.9186970 -  3.9206448
     "00100010010001000100010010001000",  --  3.9207076 -  3.9226554
     "10001001000100010001001000100010",  --  3.9227183 -  3.9246660
     "00100100010001000100100010001000",  --  3.9247289 -  3.9266767
     "10001001000100010001001000100010",  --  3.9267395 -  3.9286873
     "00100010010001000100010010001000",  --  3.9287501 -  3.9306979
     "10001000100100010001000100100010",  --  3.9307607 -  3.9327085
     "00100010001001000100010001000100",  --  3.9327713 -  3.9347191
     "10001000100010001001000100010001",  --  3.9347820 -  3.9367298
     "00010010001000100010001001000100",  --  3.9367926 -  3.9387404
     "01000100010010001000100010001000",  --  3.9388032 -  3.9407510
     "10010001000100010001001000100010",  --  3.9408138 -  3.9427616
     "00100010001001000100010001000100",  --  3.9428244 -  3.9447722
     "01001000100010001000100010010001",  --  3.9448351 -  3.9467829
     "00010001000100010010001000100010",  --  3.9468457 -  3.9487935
     "00100010010001000100010001000100",  --  3.9488563 -  3.9508041
     "01001000100010001000100010001001",  --  3.9508669 -  3.9528147
     "00010001000100010001000100100010",  --  3.9528775 -  3.9548253
     "00100010001000100010010001000100",  --  3.9548882 -  3.9568359
     "01000100010001000100100010001000",  --  3.9568988 -  3.9588466
     "10001000100010001001000100010001",  --  3.9589094 -  3.9608572
     "00010001000100010001001000100010",  --  3.9609200 -  3.9628678
     "00100010001000100010001001000100",  --  3.9629306 -  3.9648784
     "01000100010001000100010001000100",  --  3.9649413 -  3.9668890
     "10001000100010001000100010001000",  --  3.9669519 -  3.9688997
     "10001000100100010001000100010001",  --  3.9689625 -  3.9709103
     "00010001000100010001000100010010",  --  3.9709731 -  3.9729209
     "00100010001000100010001000100010",  --  3.9729837 -  3.9749315
     "00100010001000100010001001000100",  --  3.9749944 -  3.9769421
     "01000100010001000100010001000100",  --  3.9770050 -  3.9789528
     "01000100010001000100010001000100",  --  3.9790156 -  3.9809634
     "10001000100010001000100010001000",  --  3.9810262 -  3.9829740
     "10001000100010001000100010001000",  --  3.9830368 -  3.9849846
     "10001000100010001000100010001000",  --  3.9850474 -  3.9869952
     "10001000100010001000100100010001",  --  3.9870581 -  3.9890059
     "00010001000100010001000100010001",  --  3.9890687 -  3.9910165
     "00010001000100010001000100010001",  --  3.9910793 -  3.9930271
     "00010001000100010001000100010001",  --  3.9930899 -  3.9950377
     "00010001000100010001000100010001",  --  3.9951005 -  3.9970483
     "00010001000100010001000100010001",  --  3.9971112 -  3.9990590
     "00010001000100001000100010001000",  --  3.9991218 -  4.0010696
     "10001000100010001000100010001000",  --  4.0011324 -  4.0030802
     "10001000100010001000100010001000",  --  4.0031430 -  4.0050908
     "10001000100010001000100010001000",  --  4.0051536 -  4.0071014
     "10001000010001000100010001000100",  --  4.0071643 -  4.0091120
     "01000100010001000100010001000100",  --  4.0091749 -  4.0111227
     "01000100010001000010001000100010",  --  4.0111855 -  4.0131333
     "00100010001000100010001000100010",  --  4.0131961 -  4.0151439
     "00100010001000010001000100010001",  --  4.0152067 -  4.0171545
     "00010001000100010001000100010000",  --  4.0172174 -  4.0191651
     "10001000100010001000100010001000",  --  4.0192280 -  4.0211758
     "10001000100001000100010001000100",  --  4.0212386 -  4.0231864
     "01000100010001000100001000100010",  --  4.0232492 -  4.0251970
     "00100010001000100010001000010001",  --  4.0252598 -  4.0272076
     "00010001000100010001000100001000",  --  4.0272705 -  4.0292182
     "10001000100010001000100010000100",  --  4.0292811 -  4.0312289
     "01000100010001000100010001000010",  --  4.0312917 -  4.0332395
     "00100010001000100010001000010001",  --  4.0333023 -  4.0352501
     "00010001000100010001000010001000",  --  4.0353129 -  4.0372607
     "10001000100010000100010001000100",  --  4.0373236 -  4.0392713
     "01000100001000100010001000100010",  --  4.0393342 -  4.0412820
     "00100001000100010001000100001000",  --  4.0413448 -  4.0432926
     "10001000100010001000010001000100",  --  4.0433554 -  4.0453032
     "01000100010000100010001000100010",  --  4.0453660 -  4.0473138
     "00010001000100010001000010001000",  --  4.0473766 -  4.0493244
     "10001000100001000100010001000100",  --  4.0493873 -  4.0513351
     "00100010001000100010000100010001",  --  4.0513979 -  4.0533457
     "00010001000010001000100010001000",  --  4.0534085 -  4.0553563
     "01000100010001000010001000100010",  --  4.0554191 -  4.0573669
     "00100001000100010001000010001000",  --  4.0574297 -  4.0593775
     "10001000010001000100010001000010",  --  4.0594404 -  4.0613882
     "00100010001000010001000100010000",  --  4.0614510 -  4.0633988
     "10001000100010000100010001000100",  --  4.0634616 -  4.0654094
     "00100010001000100001000100010001",  --  4.0654722 -  4.0674200
     "00001000100010000100010001000100",  --  4.0674828 -  4.0694306
     "00100010001000100001000100010001",  --  4.0694935 -  4.0714412
     "00001000100010000100010001000100",  --  4.0715041 -  4.0734519
     "00100010001000010001000100010000",  --  4.0735147 -  4.0754625
     "10001000100001000100010001000010",  --  4.0755253 -  4.0774731
     "00100010000100010001000010001000",  --  4.0775359 -  4.0794837
     "10001000010001000100001000100010",  --  4.0795466 -  4.0814943
     "00010001000100001000100010000100",  --  4.0815572 -  4.0835050
     "01000100001000100010001000010001",  --  4.0835678 -  4.0855156
     "00010000100010001000010001000100",  --  4.0855784 -  4.0875262
     "00100010001000010001000100001000",  --  4.0875890 -  4.0895368
     "10001000010001000010001000100001",  --  4.0895997 -  4.0915474
     "00010001000010001000100001000100",  --  4.0916103 -  4.0935581
     "01000010001000100001000100001000",  --  4.0936209 -  4.0955687
     "10001000010001000100001000100010",  --  4.0956315 -  4.0975793
     "00010001000010001000100001000100",  --  4.0976421 -  4.0995899
     "01000010001000010001000100001000",  --  4.0996527 -  4.1016005
     "10000100010001000010001000100001",  --  4.1016634 -  4.1036112
     "00010000100010001000010001000010",  --  4.1036740 -  4.1056218
     "00100010000100010000100010001000",  --  4.1056846 -  4.1076324
     "01000100001000100001000100010000",  --  4.1076952 -  4.1096430
     "10001000010001000100001000100001",  --  4.1097058 -  4.1116536
     "00010000100010001000010001000010",  --  4.1117165 -  4.1136643
     "00100001000100010000100010000100",  --  4.1137271 -  4.1156749
     "01000010001000100001000100001000",  --  4.1157377 -  4.1176855
     "10000100010000100010001000010001",  --  4.1177483 -  4.1196961
     "00001000100001000100001000100001",  --  4.1197589 -  4.1217067
     "00010001000010001000010001000010",  --  4.1217696 -  4.1237173
     "00100001000100001000100001000100",  --  4.1237802 -  4.1257280
     "00100010001000010001000010001000",  --  4.1257908 -  4.1277386
     "01000100001000100001000100001000",  --  4.1278014 -  4.1297492
     "10000100010000100010000100010000",  --  4.1298120 -  4.1317598
     "10001000010001000010001000010001",  --  4.1318227 -  4.1337704
     "00001000100001000100001000100001",  --  4.1338333 -  4.1357811
     "00010000100010000100010000100010",  --  4.1358439 -  4.1377917
     "00010001000010001000010000100010",  --  4.1378545 -  4.1398023
     "00010001000010001000010001000010",  --  4.1398651 -  4.1418129
     "00100001000100001000100001000100",  --  4.1418758 -  4.1438235
     "00100001000100001000100001000100",  --  4.1438864 -  4.1458342
     "00100010000100010000100001000100",  --  4.1458970 -  4.1478448
     "00100010000100010000100001000100",  --  4.1479076 -  4.1498554
     "00100010000100010000100010000100",  --  4.1499182 -  4.1518660
     "00100010000100010000100010000100",  --  4.1519289 -  4.1538766
     "00100010000100010000100001000100",  --  4.1539395 -  4.1558873
     "00100010000100010000100001000100",  --  4.1559501 -  4.1578979
     "00100010000100001000100001000100",  --  4.1579607 -  4.1599085
     "00100001000100001000100001000010",  --  4.1599713 -  4.1619191
     "00100001000100001000010001000010",  --  4.1619819 -  4.1639297
     "00010001000010001000010000100010",  --  4.1639926 -  4.1659404
     "00010001000010000100010000100001",  --  4.1660032 -  4.1679510
     "00010000100010000100001000100001",  --  4.1680138 -  4.1699616
     "00001000100001000010001000010000",  --  4.1700244 -  4.1719722
     "10001000010001000010000100010000",  --  4.1720350 -  4.1739828
     "10000100010000100001000100001000",  --  4.1740457 -  4.1759935
     "01000100001000010001000010000100",  --  4.1760563 -  4.1780041
     "01000010000100010000100001000100",  --  4.1780669 -  4.1800147
     "00100001000100001000010001000010",  --  4.1800775 -  4.1820253
     "00010001000010000100010000100001",  --  4.1820881 -  4.1840359
     "00001000100001000010001000010000",  --  4.1840988 -  4.1860465
     "10001000010000100010000100001000",  --  4.1861094 -  4.1880572
     "01000100001000010001000010000100",  --  4.1881200 -  4.1900678
     "00100010000100001000100001000010",  --  4.1901306 -  4.1920784
     "00010001000010000100010000100001",  --  4.1921412 -  4.1940890
     "00001000100001000010000100010000",  --  4.1941519 -  4.1960996
     "10000100010000100001000010001000",  --  4.1961625 -  4.1981103
     "01000010000100010000100001000010",  --  4.1981731 -  4.2001209
     "00100001000010000100010000100001",  --  4.2001837 -  4.2021315
     "00001000100001000010000100010000",  --  4.2021943 -  4.2041421
     "10000100001000100001000010000100",  --  4.2042050 -  4.2061527
     "00100010000100001000010001000010",  --  4.2062156 -  4.2081634
     "00010000100001000100001000010000",  --  4.2082262 -  4.2101740
     "10001000010000100001000010001000",  --  4.2102368 -  4.2121846
     "01000010000100001000100001000010",  --  4.2122474 -  4.2141952
     "00010000100010000100001000010000",  --  4.2142580 -  4.2162058
     "10001000010000100001000010001000",  --  4.2162687 -  4.2182165
     "01000010000100001000010001000010",  --  4.2182793 -  4.2202271
     "00010000100001000100001000010000",  --  4.2202899 -  4.2222377
     "10000100001000100001000010000100",  --  4.2223005 -  4.2242483
     "00100001000100001000010000100001",  --  4.2243111 -  4.2262589
     "00001000010001000010000100001000",  --  4.2263218 -  4.2282696
     "01000010001000010000100001000010",  --  4.2283324 -  4.2302802
     "00010000100010000100001000010000",  --  4.2303430 -  4.2322908
     "10000100001000010001000010000100",  --  4.2323536 -  4.2343014
     "00100001000010000100010000100001",  --  4.2343642 -  4.2363120
     "00001000010000100001000010000100",  --  4.2363749 -  4.2383226
     "01000010000100001000010000100001",  --  4.2383855 -  4.2403333
     "00001000010001000010000100001000",  --  4.2403961 -  4.2423439
     "01000010000100001000010000100010",  --  4.2424067 -  4.2443545
     "00010000100001000010000100001000",  --  4.2444173 -  4.2463651
     "01000010000100001000010001000010",  --  4.2464280 -  4.2483757
     "00010000100001000010000100001000",  --  4.2484386 -  4.2503864
     "01000010000100001000010000100010",  --  4.2504492 -  4.2523970
     "00010000100001000010000100001000",  --  4.2524598 -  4.2544076
     "01000010000100001000010000100001",  --  4.2544704 -  4.2564182
     "00001000010000100001000010000100",  --  4.2564811 -  4.2584288
     "01000010000100001000010000100001",  --  4.2584917 -  4.2604395
     "00001000010000100001000010000100",  --  4.2605023 -  4.2624501
     "00100001000010000100001000010000",  --  4.2625129 -  4.2644607
     "10000100001000010000100001000010",  --  4.2645235 -  4.2664713
     "00010000100001000010000100001000",  --  4.2665342 -  4.2684819
     "01000010000100001000010000100001",  --  4.2685448 -  4.2704926
     "00001000010000100001000010000100",  --  4.2705554 -  4.2725032
     "00100001000010000100001000010000",  --  4.2725660 -  4.2745138
     "10000100001000010000100001000010",  --  4.2745766 -  4.2765244
     "00010000100001000010000100001000",  --  4.2765872 -  4.2785350
     "01000010000100001000010000100001",  --  4.2785979 -  4.2805457
     "00001000001000010000100001000010",  --  4.2806085 -  4.2825563
     "00010000100001000010000100001000",  --  4.2826191 -  4.2845669
     "01000010000100001000010000100001",  --  4.2846297 -  4.2865775
     "00001000010000010000100001000010",  --  4.2866403 -  4.2885881
     "00010000100001000010000100001000",  --  4.2886510 -  4.2905988
     "01000010000100001000001000010000",  --  4.2906616 -  4.2926094
     "10000100001000010000100001000010",  --  4.2926722 -  4.2946200
     "00010000100001000001000010000100",  --  4.2946828 -  4.2966306
     "00100001000010000100001000010000",  --  4.2966934 -  4.2986412
     "10000010000100001000010000100001",  --  4.2987041 -  4.3006518
     "00001000010000100000100001000010",  --  4.3007147 -  4.3026625
     "00010000100001000010000100001000",  --  4.3027253 -  4.3046731
     "00100001000010000100001000010000",  --  4.3047359 -  4.3066837
     "10000100000100001000010000100001",  --  4.3067465 -  4.3086943
     "00001000010000010000100001000010",  --  4.3087572 -  4.3107049
     "00010000100001000001000010000100",  --  4.3107678 -  4.3127156
     "00100001000010000100000100001000",  --  4.3127784 -  4.3147262
     "01000010000100001000001000010000",  --  4.3147890 -  4.3167368
     "10000100001000010000010000100001",  --  4.3167996 -  4.3187474
     "00001000010000100000100001000010",  --  4.3188103 -  4.3207580
     "00010000100001000001000010000100",  --  4.3208209 -  4.3227687
     "00100001000001000010000100001000",  --  4.3228315 -  4.3247793
     "01000001000010000100001000010000",  --  4.3248421 -  4.3267899
     "10000010000100001000010000100000",  --  4.3268527 -  4.3288005
     "10000100001000010000010000100001",  --  4.3288633 -  4.3308111
     "00001000010000010000100001000010",  --  4.3308740 -  4.3328218
     "00010000010000100001000010000010",  --  4.3328846 -  4.3348324
     "00010000100001000010000010000100",  --  4.3348952 -  4.3368430
     "00100001000001000010000100001000",  --  4.3369058 -  4.3388536
     "00100001000010000100000100001000",  --  4.3389164 -  4.3408642
     "01000010000010000100001000010000",  --  4.3409271 -  4.3428749
     "01000010000100001000001000010000",  --  4.3429377 -  4.3448855
     "10000100000100001000010000100000",  --  4.3449483 -  4.3468961
     "10000100001000010000010000100001",  --  4.3469589 -  4.3489067
     "00000100001000010000100000100001",  --  4.3489695 -  4.3509173
     "00001000010000010000100001000001",  --  4.3509802 -  4.3529279
     "00001000010000100000100001000010",  --  4.3529908 -  4.3549386
     "00001000010000100001000001000010",  --  4.3550014 -  4.3569492
     "00010000010000100001000001000010",  --  4.3570120 -  4.3589598
     "00010000100000100001000010000010",  --  4.3590226 -  4.3609704
     "00010000100000100001000010000010",  --  4.3610333 -  4.3629810
     "00010000100000100001000010000010",  --  4.3630439 -  4.3649917
     "00010000100000100001000010000100",  --  4.3650545 -  4.3670023
     "00010000100001000001000010000100",  --  4.3670651 -  4.3690129
     "00010000100000100001000010000010",  --  4.3690757 -  4.3710235
     "00010000100000100001000010000010",  --  4.3710864 -  4.3730341
     "00010000100000100001000010000010",  --  4.3730970 -  4.3750448
     "00010000100000100001000001000010",  --  4.3751076 -  4.3770554
     "00010000010000100001000001000010",  --  4.3771182 -  4.3790660
     "00010000010000100000100001000010",  --  4.3791288 -  4.3810766
     "00001000010000100000100001000001",  --  4.3811395 -  4.3830872
     "00001000010000010000100001000001",  --  4.3831501 -  4.3850979
     "00001000001000010000100000100001",  --  4.3851607 -  4.3871085
     "00000100001000010000010000100000",  --  4.3871713 -  4.3891191
     "10000100001000001000010000010000",  --  4.3891819 -  4.3911297
     "10000100000100001000001000010000",  --  4.3911925 -  4.3931403
     "10000010000100000100001000001000",  --  4.3932032 -  4.3951510
     "01000010000010000100000100001000",  --  4.3952138 -  4.3971616
     "01000001000010000010000100000100",  --  4.3972244 -  4.3991722
     "00100001000001000010000010000100",  --  4.3992350 -  4.4011828
     "00010000100000100001000010000010",  --  4.4012456 -  4.4031934
     "00010000010000100000100001000010",  --  4.4032563 -  4.4052041
     "00001000010000010000100000100001",  --  4.4052669 -  4.4072147
     "00000100001000001000010000100000",  --  4.4072775 -  4.4092253
     "10000100000100001000001000010000",  --  4.4092881 -  4.4112359
     "01000010000010000100000100001000",  --  4.4112987 -  4.4132465
     "00100001000010000010000100000100",  --  4.4133094 -  4.4152571
     "00100000100001000001000010000010",  --  4.4153200 -  4.4172678
     "00010000010000100000100001000001",  --  4.4173306 -  4.4192784
     "00001000001000010000010000100000",  --  4.4193412 -  4.4212890
     "10000100000100001000001000010000",  --  4.4213518 -  4.4232996
     "01000010000010000100000100001000",  --  4.4233625 -  4.4253102
     "00100001000001000010000010000100",  --  4.4253731 -  4.4273209
     "00010000100000100001000001000010",  --  4.4273837 -  4.4293315
     "00001000010000010000100000100001",  --  4.4293943 -  4.4313421
     "00000100000100001000001000010000",  --  4.4314049 -  4.4333527
     "01000010000010000100000100001000",  --  4.4334156 -  4.4353633
     "00100001000001000010000010000010",  --  4.4354262 -  4.4373740
     "00010000010000100000100001000001",  --  4.4374368 -  4.4393846
     "00001000001000010000010000010000",  --  4.4394474 -  4.4413952
     "10000010000100000100001000001000",  --  4.4414580 -  4.4434058
     "01000001000001000010000010000100",  --  4.4434686 -  4.4454164
     "00010000100000100001000001000001",  --  4.4454793 -  4.4474271
     "00001000001000010000010000100000",  --  4.4474899 -  4.4494377
     "10000010000100000100001000001000",  --  4.4495005 -  4.4514483
     "01000001000001000010000010000100",  --  4.4515111 -  4.4534589
     "00010000010000100000100001000001",  --  4.4535217 -  4.4554695
     "00001000001000001000010000010000",  --  4.4555324 -  4.4574802
     "10000010000010000100000100001000",  --  4.4575430 -  4.4594908
     "00100000100001000001000010000010",  --  4.4595536 -  4.4615014
     "00001000010000010000100000100000",  --  4.4615642 -  4.4635120
     "10000100000100000100001000001000",  --  4.4635748 -  4.4655226
     "01000001000001000010000010000100",  --  4.4655855 -  4.4675332
     "00010000010000100000100000100001",  --  4.4675961 -  4.4695439
     "00000100001000001000001000010000",  --  4.4696067 -  4.4715545
     "01000001000010000010000010000100",  --  4.4716173 -  4.4735651
     "00010000100000100000100001000001",  --  4.4736279 -  4.4755757
     "00000100001000001000001000010000",  --  4.4756386 -  4.4775863
     "01000001000010000010000100000100",  --  4.4776492 -  4.4795970
     "00010000100000100000100001000001",  --  4.4796598 -  4.4816076
     "00000100001000001000001000010000",  --  4.4816704 -  4.4836182
     "01000001000010000010000010000100",  --  4.4836810 -  4.4856288
     "00010000010000100000100000100001",  --  4.4856917 -  4.4876394
     "00000100000100001000001000001000",  --  4.4877023 -  4.4896501
     "01000001000001000010000010000010",  --  4.4897129 -  4.4916607
     "00010000010000010000100000100000",  --  4.4917235 -  4.4936713
     "10000010000100000100000100001000",  --  4.4937341 -  4.4956819
     "00100000100001000001000001000010",  --  4.4957448 -  4.4976925
     "00001000001000010000010000010000",  --  4.4977554 -  4.4997032
     "01000010000010000010000100000100",  --  4.4997660 -  4.5017138
     "00010000100000100000100000100001",  --  4.5017766 -  4.5037244
     "00000100000100001000001000001000",  --  4.5037872 -  4.5057350
     "00100001000001000001000010000010",  --  4.5057978 -  4.5077456
     "00001000001000010000010000010000",  --  4.5078085 -  4.5097563
     "10000010000010000010000100000100",  --  4.5098191 -  4.5117669
     "00010000010000100000100000100001",  --  4.5118297 -  4.5137775
     "00000100000100000100001000001000",  --  4.5138403 -  4.5157881
     "00100000100001000001000001000001",  --  4.5158509 -  4.5177987
     "00001000001000001000010000010000",  --  4.5178616 -  4.5198094
     "01000001000010000010000010000010",  --  4.5198722 -  4.5218200
     "00010000010000010000010000100000",  --  4.5218828 -  4.5238306
     "10000010000010000100000100000100",  --  4.5238934 -  4.5258412
     "00010000100000100000100000100001",  --  4.5259040 -  4.5278518
     "00000100000100000100000100001000",  --  4.5279147 -  4.5298624
     "00100000100000100001000001000001",  --  4.5299253 -  4.5318731
     "00000100001000001000001000001000",  --  4.5319359 -  4.5338837
     "01000001000001000001000001000010",  --  4.5339465 -  4.5358943
     "00001000001000001000010000010000",  --  4.5359571 -  4.5379049
     "01000001000001000010000010000010",  --  4.5379678 -  4.5399155
     "00001000010000010000010000010000",  --  4.5399784 -  4.5419262
     "01000010000010000010000010000010",  --  4.5419890 -  4.5439368
     "00010000010000010000010000010000",  --  4.5439996 -  4.5459474
     "10000010000010000010000010000100",  --  4.5460102 -  4.5479580
     "00010000010000010000010000100000",  --  4.5480209 -  4.5499686
     "10000010000010000010000100000100",  --  4.5500315 -  4.5519793
     "00010000010000010000100000100000",  --  4.5520421 -  4.5539899
     "10000010000010000100000100000100",  --  4.5540527 -  4.5560005
     "00010000010000100000100000100000",  --  4.5560633 -  4.5580111
     "10000010000010000100000100000100",  --  4.5580739 -  4.5600217
     "00010000010000100000100000100000",  --  4.5600846 -  4.5620324
     "10000010000010000100000100000100",  --  4.5620952 -  4.5640430
     "00010000010000010000100000100000",  --  4.5641058 -  4.5660536
     "10000010000010000100000100000100",  --  4.5661164 -  4.5680642
     "00010000010000010000100000100000",  --  4.5681270 -  4.5700748
     "10000010000010000010000010000100",  --  4.5701377 -  4.5720855
     "00010000010000010000010000010000",  --  4.5721483 -  4.5740961
     "10000010000010000010000010000010",  --  4.5741589 -  4.5761067
     "00010000010000010000010000010000",  --  4.5761695 -  4.5781173
     "01000001000010000010000010000010",  --  4.5781801 -  4.5801279
     "00001000001000010000010000010000",  --  4.5801908 -  4.5821385
     "01000001000001000001000010000010",  --  4.5822014 -  4.5841492
     "00001000001000001000001000001000",  --  4.5842120 -  4.5861598
     "01000001000001000001000001000001",  --  4.5862226 -  4.5881704
     "00000100000100001000001000001000",  --  4.5882332 -  4.5901810
     "00100000100000100000100001000001",  --  4.5902439 -  4.5921916
     "00000100000100000100000100000100",  --  4.5922545 -  4.5942023
     "00010000100000100000100000100000",  --  4.5942651 -  4.5962129
     "10000010000010000010000100000100",  --  4.5962757 -  4.5982235
     "00010000010000010000010000010000",  --  4.5982863 -  4.6002341
     "01000010000010000010000010000010",  --  4.6002970 -  4.6022447
     "00001000001000001000010000010000",  --  4.6023076 -  4.6042554
     "01000001000001000001000001000001",  --  4.6043182 -  4.6062660
     "00000100001000001000001000001000",  --  4.6063288 -  4.6082766
     "00100000100000100000100000100001",  --  4.6083394 -  4.6102872
     "00000100000100000100000100000100",  --  4.6103501 -  4.6122978
     "00010000010000010000010000100000",  --  4.6123607 -  4.6143085
     "10000010000010000010000010000010",  --  4.6143713 -  4.6163191
     "00001000001000010000010000010000",  --  4.6163819 -  4.6183297
     "01000001000001000001000001000001",  --  4.6183925 -  4.6203403
     "00000100001000001000001000001000",  --  4.6204031 -  4.6223509
     "00100000100000100000100000100000",  --  4.6224138 -  4.6243616
     "10000010000100000100000100000100",  --  4.6244244 -  4.6263722
     "00010000010000010000010000010000",  --  4.6264350 -  4.6283828
     "01000001000010000010000010000010",  --  4.6284456 -  4.6303934
     "00001000001000001000001000001000",  --  4.6304562 -  4.6324040
     "00100000100000100001000001000001",  --  4.6324669 -  4.6344147
     "00000100000100000100000100000100",  --  4.6344775 -  4.6364253
     "00010000010000010000010000100000",  --  4.6364881 -  4.6384359
     "10000010000010000010000010000010",  --  4.6384987 -  4.6404465
     "00001000001000001000001000001000",  --  4.6405093 -  4.6424571
     "00100001000001000001000001000001",  --  4.6425200 -  4.6444677
     "00000100000100000100000100000100",  --  4.6445306 -  4.6464784
     "00010000010000010000100000100000",  --  4.6465412 -  4.6484890
     "10000010000010000010000010000010",  --  4.6485518 -  4.6504996
     "00001000001000001000001000001000",  --  4.6505624 -  4.6525102
     "00100000100001000001000001000001",  --  4.6525731 -  4.6545208
     "00000100000100000100000100000100",  --  4.6545837 -  4.6565315
     "00010000010000010000010000010000",  --  4.6565943 -  4.6585421
     "01000010000010000010000010000010",  --  4.6586049 -  4.6605527
     "00001000001000001000001000001000",  --  4.6606155 -  4.6625633
     "00100000100000100000100000100000",  --  4.6626262 -  4.6645739
     "10000100000100000100000100000100",  --  4.6646368 -  4.6665846
     "00010000010000010000010000010000",  --  4.6666474 -  4.6685952
     "01000001000001000001000001000001",  --  4.6686580 -  4.6706058
     "00001000001000001000001000001000",  --  4.6706686 -  4.6726164
     "00100000100000100000100000100000",  --  4.6726792 -  4.6746270
     "10000010000010000010000010000010",  --  4.6746899 -  4.6766377
     "00001000001000010000010000010000",  --  4.6767005 -  4.6786483
     "01000001000001000001000001000001",  --  4.6787111 -  4.6806589
     "00000100000100000100000100000100",  --  4.6807217 -  4.6826695
     "00010000010000010000010000010000",  --  4.6827323 -  4.6846801
     "10000010000010000010000010000010",  --  4.6847430 -  4.6866908
     "00001000001000001000001000001000",  --  4.6867536 -  4.6887014
     "00100000100000100000100000100000",  --  4.6887642 -  4.6907120
     "10000010000010000100000100000100",  --  4.6907748 -  4.6927226
     "00010000010000010000010000010000",  --  4.6927854 -  4.6947332
     "01000001000001000001000001000001",  --  4.6947961 -  4.6967438
     "00000100000100000100000100000100",  --  4.6968067 -  4.6987545
     "00010000010000100000100000100000",  --  4.6988173 -  4.7007651
     "10000010000010000010000010000010",  --  4.7008279 -  4.7027757
     "00001000001000001000001000001000",  --  4.7028385 -  4.7047863
     "00100000100000100000100000100000",  --  4.7048492 -  4.7067969
     "10000010000100000100000100000100",  --  4.7068598 -  4.7088076
     "00010000010000010000010000010000",  --  4.7088704 -  4.7108182
     "01000001000001000001000001000001",  --  4.7108810 -  4.7128288
     "00000100000100000100000100000100",  --  4.7128916 -  4.7148394
     "00100000100000100000100000100000",  --  4.7149023 -  4.7168500
     "10000010000010000010000010000010",  --  4.7169129 -  4.7188607
     "00001000001000001000001000001000",  --  4.7189235 -  4.7208713
     "00100000100000100000100000100001",  --  4.7209341 -  4.7228819
     "00000100000100000100000100000100",  --  4.7229447 -  4.7248925
     "00010000010000010000010000010000",  --  4.7249554 -  4.7269031
     "01000001000001000001000001000001",  --  4.7269660 -  4.7289138
     "00000100000100000100000100001000",  --  4.7289766 -  4.7309244
     "00100000100000100000100000100000",  --  4.7309872 -  4.7329350
     "10000010000010000010000010000010",  --  4.7329978 -  4.7349456
     "00001000001000001000001000001000",  --  4.7350084 -  4.7369562
     "00100000100000100001000001000001",  --  4.7370191 -  4.7389669
     "00000100000100000100000100000100",  --  4.7390297 -  4.7409775
     "00010000010000010000010000010000",  --  4.7410403 -  4.7429881
     "01000001000001000001000001000001",  --  4.7430509 -  4.7449987
     "00001000001000001000001000001000",  --  4.7450615 -  4.7470093
     "00100000100000100000100000100000",  --  4.7470722 -  4.7490200
     "10000010000010000010000010000010",  --  4.7490828 -  4.7510306
     "00001000001000010000010000010000",  --  4.7510934 -  4.7530412
     "01000001000001000001000001000001",  --  4.7531040 -  4.7550518
     "00000100000100000100000100000100",  --  4.7551146 -  4.7570624
     "00010000010000010000100000100000",  --  4.7571253 -  4.7590730
     "10000010000010000010000010000010",  --  4.7591359 -  4.7610837
     "00001000001000001000001000001000",  --  4.7611465 -  4.7630943
     "00100000100000100001000001000001",  --  4.7631571 -  4.7651049
     "00000100000100000100000100000100",  --  4.7651677 -  4.7671155
     "00010000010000010000010000010000",  --  4.7671784 -  4.7691261
     "01000001000010000010000010000010",  --  4.7691890 -  4.7711368
     "00001000001000001000001000001000",  --  4.7711996 -  4.7731474
     "00100000100000100000100000100000",  --  4.7732102 -  4.7751580
     "10000100000100000100000100000100",  --  4.7752208 -  4.7771686
     "00010000010000010000010000010000",  --  4.7772315 -  4.7791792
     "01000001000001000001000010000010",  --  4.7792421 -  4.7811899
     "00001000001000001000001000001000",  --  4.7812527 -  4.7832005
     "00100000100000100000100000100000",  --  4.7832633 -  4.7852111
     "10000100000100000100000100000100",  --  4.7852739 -  4.7872217
     "00010000010000010000010000010000",  --  4.7872845 -  4.7892323
     "01000001000010000010000010000010",  --  4.7892952 -  4.7912430
     "00001000001000001000001000001000",  --  4.7913058 -  4.7932536
     "00100000100000100001000001000001",  --  4.7933164 -  4.7952642
     "00000100000100000100000100000100",  --  4.7953270 -  4.7972748
     "00010000010000010000100000100000",  --  4.7973376 -  4.7992854
     "10000010000010000010000010000010",  --  4.7993483 -  4.8012961
     "00001000001000001000010000010000",  --  4.8013589 -  4.8033067
     "01000001000001000001000001000001",  --  4.8033695 -  4.8053173
     "00000100000100001000001000001000",  --  4.8053801 -  4.8073279
     "00100000100000100000100000100000",  --  4.8073907 -  4.8093385
     "10000010000100000100000100000100",  --  4.8094014 -  4.8113491
     "00010000010000010000010000010000",  --  4.8114120 -  4.8133598
     "01000010000010000010000010000010",  --  4.8134226 -  4.8153704
     "00001000001000001000001000010000",  --  4.8154332 -  4.8173810
     "01000001000001000001000001000001",  --  4.8174438 -  4.8193916
     "00000100000100001000001000001000",  --  4.8194545 -  4.8214022
     "00100000100000100000100000100001",  --  4.8214651 -  4.8234129
     "00000100000100000100000100000100",  --  4.8234757 -  4.8254235
     "00010000010000010000100000100000",  --  4.8254863 -  4.8274341
     "10000010000010000010000010000010",  --  4.8274969 -  4.8294447
     "00010000010000010000010000010000",  --  4.8295076 -  4.8314553
     "01000001000010000010000010000010",  --  4.8315182 -  4.8334660
     "00001000001000001000001000010000",  --  4.8335288 -  4.8354766
     "01000001000001000001000001000001",  --  4.8355394 -  4.8374872
     "00001000001000001000001000001000",  --  4.8375500 -  4.8394978
     "00100000100001000001000001000001",  --  4.8395607 -  4.8415084
     "00000100000100000100001000001000",  --  4.8415713 -  4.8435191
     "00100000100000100000100000100001",  --  4.8435819 -  4.8455297
     "00000100000100000100000100000100",  --  4.8455925 -  4.8475403
     "00010000100000100000100000100000",  --  4.8476031 -  4.8495509
     "10000010000100000100000100000100",  --  4.8496137 -  4.8515615
     "00010000010000100000100000100000",  --  4.8516244 -  4.8535722
     "10000010000010000100000100000100",  --  4.8536350 -  4.8555828
     "00010000010000010000010000100000",  --  4.8556456 -  4.8575934
     "10000010000010000010000100000100",  --  4.8576562 -  4.8596040
     "00010000010000010000010000100000",  --  4.8596668 -  4.8616146
     "10000010000010000010000010000100",  --  4.8616775 -  4.8636253
     "00010000010000010000010000100000",  --  4.8636881 -  4.8656359
     "10000010000010000010000010000100",  --  4.8656987 -  4.8676465
     "00010000010000010000010000100000",  --  4.8677093 -  4.8696571
     "10000010000010000010000100000100",  --  4.8697199 -  4.8716677
     "00010000010000010000010000100000",  --  4.8717306 -  4.8736783
     "10000010000010000010000100000100",  --  4.8737412 -  4.8756890
     "00010000010000010000100000100000",  --  4.8757518 -  4.8776996
     "10000010000010000100000100000100",  --  4.8777624 -  4.8797102
     "00010000100000100000100000100000",  --  4.8797730 -  4.8817208
     "10000100000100000100000100000100",  --  4.8817837 -  4.8837314
     "00100000100000100000100000100001",  --  4.8837943 -  4.8857421
     "00000100000100000100001000001000",  --  4.8858049 -  4.8877527
     "00100000100000100001000001000001",  --  4.8878155 -  4.8897633
     "00000100001000001000001000001000",  --  4.8898261 -  4.8917739
     "01000001000001000001000001000010",  --  4.8918368 -  4.8937845
     "00001000001000001000010000010000",  --  4.8938474 -  4.8957952
     "01000001000010000010000010000010",  --  4.8958580 -  4.8978058
     "00010000010000010000010000100000",  --  4.8978686 -  4.8998164
     "10000010000010000100000100000100",  --  4.8998792 -  4.9018270
     "00010000100000100000100000100001",  --  4.9018898 -  4.9038376
     "00000100000100000100001000001000",  --  4.9039005 -  4.9058483
     "00100000100001000001000001000001",  --  4.9059111 -  4.9078589
     "00001000001000001000001000010000",  --  4.9079217 -  4.9098695
     "01000001000010000010000010000010",  --  4.9099323 -  4.9118801
     "00010000010000010000010000100000",  --  4.9119429 -  4.9138907
     "10000010000100000100000100000100",  --  4.9139536 -  4.9159014
     "00100000100000100001000001000001",  --  4.9159642 -  4.9179120
     "00000100001000001000001000010000",  --  4.9179748 -  4.9199226
     "01000001000001000010000010000010",  --  4.9199854 -  4.9219332
     "00010000010000010000010000100000",  --  4.9219960 -  4.9239438
     "10000010000100000100000100001000",  --  4.9240067 -  4.9259544
     "00100000100000100001000001000001",  --  4.9260173 -  4.9279651
     "00001000001000001000010000010000",  --  4.9280279 -  4.9299757
     "01000010000010000010000100000100",  --  4.9300385 -  4.9319863
     "00010000010000100000100000100001",  --  4.9320491 -  4.9339969
     "00000100000100001000001000001000",  --  4.9340598 -  4.9360075
     "01000001000001000010000010000010",  --  4.9360704 -  4.9380182
     "00010000010000010000100000100000",  --  4.9380810 -  4.9400288
     "10000100000100000100001000001000",  --  4.9400916 -  4.9420394
     "00100001000001000001000010000010",  --  4.9421022 -  4.9440500
     "00001000010000010000010000100000",  --  4.9441129 -  4.9460606
     "10000100000100000100001000001000",  --  4.9461235 -  4.9480713
     "00100001000001000001000010000010",  --  4.9481341 -  4.9500819
     "00001000010000010000100000100000",  --  4.9501447 -  4.9520925
     "10000100000100000100001000001000",  --  4.9521553 -  4.9541031
     "00100001000001000010000010000010",  --  4.9541660 -  4.9561137
     "00010000010000010000100000100001",  --  4.9561766 -  4.9581244
     "00000100000100001000001000010000",  --  4.9581872 -  4.9601350
     "01000001000010000010000010000100",  --  4.9601978 -  4.9621456
     "00010000100000100000100001000001",  --  4.9622084 -  4.9641562
     "00001000001000001000010000010000",  --  4.9642190 -  4.9661668
     "10000010000010000100000100001000",  --  4.9662297 -  4.9681775
     "00100000100001000001000010000010",  --  4.9682403 -  4.9701881
     "00010000010000010000100000100001",  --  4.9702509 -  4.9721987
     "00000100000100001000001000010000",  --  4.9722615 -  4.9742093
     "01000010000010000010000100000100",  --  4.9742721 -  4.9762199
     "00100000100001000001000001000010",  --  4.9762828 -  4.9782306
     "00001000010000010000100000100000",  --  4.9782934 -  4.9802412
     "10000100000100001000001000010000",  --  4.9803040 -  4.9822518
     "01000010000010000010000100000100",  --  4.9823146 -  4.9842624
     "00100000100001000001000010000010",  --  4.9843252 -  4.9862730
     "00010000010000010000100000100001",  --  4.9863359 -  4.9882836
     "00000100001000001000010000010000",  --  4.9883465 -  4.9902943
     "10000010000100000100000100001000",  --  4.9903571 -  4.9923049
     "00100001000001000010000010000100",  --  4.9923677 -  4.9943155
     "00010000100000100001000001000010",  --  4.9943783 -  4.9963261
     "00001000010000010000100000100001",  --  4.9963890 -  4.9983367
     "00000100001000001000010000010000",  --  4.9983996 -  5.0003474
     "10000010000100000100001000001000",  --  5.0004102 -  5.0023580
     "01000001000010000010000100000100",  --  5.0024208 -  5.0043686
     "00100000100001000001000010000010",  --  5.0044314 -  5.0063792
     "00010000010000100000100001000001",  --  5.0064421 -  5.0083898
     "00001000001000010000010000100000",  --  5.0084527 -  5.0104005
     "10000100000100001000001000010000",  --  5.0104633 -  5.0124111
     "10000010000100000100001000001000",  --  5.0124739 -  5.0144217
     "01000001000010000010000100000100",  --  5.0144845 -  5.0164323
     "00100001000001000010000010000100",  --  5.0164951 -  5.0184429
     "00010000100000100001000001000010",  --  5.0185058 -  5.0204536
     "00010000010000100000100001000001",  --  5.0205164 -  5.0224642
     "00001000001000010000100000100001",  --  5.0225270 -  5.0244748
     "00000100001000001000010000100000",  --  5.0245376 -  5.0264854
     "10000100000100001000001000010000",  --  5.0265482 -  5.0284960
     "10000010000100000100001000001000",  --  5.0285589 -  5.0305067
     "01000010000010000100000100001000",  --  5.0305695 -  5.0325173
     "01000001000010000010000100001000",  --  5.0325801 -  5.0345279
     "00100001000001000010000100000100",  --  5.0345907 -  5.0365385
     "00100000100001000010000010000100",  --  5.0366013 -  5.0385491
     "00010000100001000001000010000010",  --  5.0386120 -  5.0405597
     "00010000100000100001000010000010",  --  5.0406226 -  5.0425704
     "00010000010000100001000001000010",  --  5.0426332 -  5.0445810
     "00010000010000100000100001000010",  --  5.0446438 -  5.0465916
     "00001000010000100000100001000010",  --  5.0466544 -  5.0486022
     "00001000010000010000100001000001",  --  5.0486651 -  5.0506128
     "00001000010000010000100001000001",  --  5.0506757 -  5.0526235
     "00001000010000010000100001000001",  --  5.0526863 -  5.0546341
     "00001000010000010000100001000001",  --  5.0546969 -  5.0566447
     "00001000010000010000100001000001",  --  5.0567075 -  5.0586553
     "00001000010000010000100001000001",  --  5.0587182 -  5.0606659
     "00001000010000010000100001000001",  --  5.0607288 -  5.0626766
     "00001000010000010000100001000010",  --  5.0627394 -  5.0646872
     "00001000010000100000100001000010",  --  5.0647500 -  5.0666978
     "00001000010000100000100001000010",  --  5.0667606 -  5.0687084
     "00010000010000100001000001000010",  --  5.0687713 -  5.0707190
     "00010000100000100001000010000010",  --  5.0707819 -  5.0727297
     "00010000100001000001000010000100",  --  5.0727925 -  5.0747403
     "00010000100001000010000010000100",  --  5.0748031 -  5.0767509
     "00100001000001000010000100001000",  --  5.0768137 -  5.0787615
     "00100001000010000010000100001000",  --  5.0788243 -  5.0807721
     "01000001000010000100001000001000",  --  5.0808350 -  5.0827828
     "01000010000100000100001000010000",  --  5.0828456 -  5.0847934
     "10000010000100001000010000100000",  --  5.0848562 -  5.0868040
     "10000100001000010000010000100001",  --  5.0868668 -  5.0888146
     "00001000001000010000100001000010",  --  5.0888774 -  5.0908252
     "00001000010000100001000001000010",  --  5.0908881 -  5.0928359
     "00010000100001000001000010000100",  --  5.0928987 -  5.0948465
     "00100001000001000010000100001000",  --  5.0949093 -  5.0968571
     "01000001000010000100001000010000",  --  5.0969199 -  5.0988677
     "01000010000100001000010000010000",  --  5.0989305 -  5.1008783
     "10000100001000010000010000100001",  --  5.1009412 -  5.1028889
     "00001000010000100000100001000010",  --  5.1029518 -  5.1048996
     "00010000100000100001000010000100",  --  5.1049624 -  5.1069102
     "00100001000001000010000100001000",  --  5.1069730 -  5.1089208
     "01000010000010000100001000010000",  --  5.1089836 -  5.1109314
     "10000100001000001000010000100001",  --  5.1109943 -  5.1129420
     "00001000010000100000100001000010",  --  5.1130049 -  5.1149527
     "00010000100001000010000010000100",  --  5.1150155 -  5.1169633
     "00100001000010000100001000001000",  --  5.1170261 -  5.1189739
     "01000010000100001000010000100001",  --  5.1190367 -  5.1209845
     "00001000001000010000100001000010",  --  5.1210474 -  5.1229951
     "00010000100001000001000010000100",  --  5.1230580 -  5.1250058
     "00100001000010000100001000010000",  --  5.1250686 -  5.1270164
     "10000010000100001000010000100001",  --  5.1270792 -  5.1290270
     "00001000010000100001000010000010",  --  5.1290898 -  5.1310376
     "00010000100001000010000100001000",  --  5.1311004 -  5.1330482
     "01000010000100001000010000100000",  --  5.1331111 -  5.1350589
     "10000100001000010000100001000010",  --  5.1351217 -  5.1370695
     "00010000100001000010000100001000",  --  5.1371323 -  5.1390801
     "01000010000100000100001000010000",  --  5.1391429 -  5.1410907
     "10000100001000010000100001000010",  --  5.1411535 -  5.1431013
     "00010000100001000010000100001000",  --  5.1431642 -  5.1451120
     "01000010000100001000010000100001",  --  5.1451748 -  5.1471226
     "00001000010000010000100001000010",  --  5.1471854 -  5.1491332
     "00010000100001000010000100001000",  --  5.1491960 -  5.1511438
     "01000010000100001000010000100001",  --  5.1512066 -  5.1531544
     "00001000010000100001000010000100",  --  5.1532173 -  5.1551650
     "00100001000010000100001000010000",  --  5.1552279 -  5.1571757
     "10000100001000010000100001000010",  --  5.1572385 -  5.1591863
     "00010000100001000010000100001000",  --  5.1592491 -  5.1611969
     "01000010000100010000100001000010",  --  5.1612597 -  5.1632075
     "00010000100001000010000100001000",  --  5.1632704 -  5.1652181
     "01000010000100001000010000100001",  --  5.1652810 -  5.1672288
     "00001000010000100001000010000100",  --  5.1672916 -  5.1692394
     "00100001000010001000010000100001",  --  5.1693022 -  5.1712500
     "00001000010000100001000010000100",  --  5.1713128 -  5.1732606
     "00100001000010000100001000010001",  --  5.1733235 -  5.1752712
     "00001000010000100001000010000100",  --  5.1753341 -  5.1772819
     "00100001000010000100001000100001",  --  5.1773447 -  5.1792925
     "00001000010000100001000010000100",  --  5.1793553 -  5.1813031
     "00100001000010001000010000100001",  --  5.1813659 -  5.1833137
     "00001000010000100001000010000100",  --  5.1833766 -  5.1853243
     "01000010000100001000010000100001",  --  5.1853872 -  5.1873350
     "00001000010001000010000100001000",  --  5.1873978 -  5.1893456
     "01000010000100001000100001000010",  --  5.1894084 -  5.1913562
     "00010000100001000010000100010000",  --  5.1914190 -  5.1933668
     "10000100001000010000100001000100",  --  5.1934296 -  5.1953774
     "00100001000010000100001000010001",  --  5.1954403 -  5.1973881
     "00001000010000100001000010001000",  --  5.1974509 -  5.1993987
     "01000010000100001000010001000010",  --  5.1994615 -  5.2014093
     "00010000100001000010001000010000",  --  5.2014721 -  5.2034199
     "10000100001000010001000010000100",  --  5.2034827 -  5.2054305
     "00100001000100001000010000100001",  --  5.2054934 -  5.2074412
     "00001000100001000010000100001000",  --  5.2075040 -  5.2094518
     "10000100001000010000100010000100",  --  5.2095146 -  5.2114624
     "00100001000010001000010000100001",  --  5.2115252 -  5.2134730
     "00001000100001000010000100010000",  --  5.2135358 -  5.2154836
     "10000100001000010001000010000100",  --  5.2155465 -  5.2174942
     "00100010000100001000010000100010",  --  5.2175571 -  5.2195049
     "00010000100001000100001000010000",  --  5.2195677 -  5.2215155
     "10001000010000100001000100001000",  --  5.2215783 -  5.2235261
     "01000010001000010000100001000100",  --  5.2235889 -  5.2255367
     "00100001000010001000010000100001",  --  5.2255996 -  5.2275473
     "00010000100001000010001000010000",  --  5.2276102 -  5.2295580
     "10001000010000100001000100001000",  --  5.2296208 -  5.2315686
     "01000010001000010000100010000100",  --  5.2316314 -  5.2335792
     "00100001000100001000010001000010",  --  5.2336420 -  5.2355898
     "00010000100010000100001000100001",  --  5.2356527 -  5.2376004
     "00001000100001000010000100010000",  --  5.2376633 -  5.2396111
     "10000100010000100001000100001000",  --  5.2396739 -  5.2416217
     "01000100001000010001000010000100",  --  5.2416845 -  5.2436323
     "00100010000100001000100001000010",  --  5.2436951 -  5.2456429
     "00100001000010001000010000100010",  --  5.2457057 -  5.2476535
     "00010000100010000100001000100001",  --  5.2477164 -  5.2496642
     "00001000100001000100001000010001",  --  5.2497270 -  5.2516748
     "00001000010001000010000100010000",  --  5.2517376 -  5.2536854
     "10000100010000100010000100001000",  --  5.2537482 -  5.2556960
     "10000100001000100001000010001000",  --  5.2557588 -  5.2577066
     "01000100001000010001000010000100",  --  5.2577695 -  5.2597173
     "01000010001000010000100010000100",  --  5.2597801 -  5.2617279
     "01000010000100010000100001000100",  --  5.2617907 -  5.2637385
     "00100010000100001000100001000100",  --  5.2638013 -  5.2657491
     "00100001000100001000100001000100",  --  5.2658119 -  5.2677597
     "00100001000100001000100001000010",  --  5.2678226 -  5.2697703
     "00100001000100001000100001000010",  --  5.2698332 -  5.2717810
     "00100001000100001000100001000010",  --  5.2718438 -  5.2737916
     "00100001000100001000100001000010",  --  5.2738544 -  5.2758022
     "00100001000100001000100001000100",  --  5.2758650 -  5.2778128
     "00100001000100001000100001000100",  --  5.2778757 -  5.2798234
     "00100010000100010000100001000100",  --  5.2798863 -  5.2818341
     "00100010000100010000100010000100",  --  5.2818969 -  5.2838447
     "01000010001000010001000010000100",  --  5.2839075 -  5.2858553
     "01000010001000010001000010001000",  --  5.2859181 -  5.2878659
     "01000100001000100001000100001000",  --  5.2879288 -  5.2898765
     "10000100010000100010000100010000",  --  5.2899394 -  5.2918872
     "10001000010001000010001000010001",  --  5.2919500 -  5.2938978
     "00001000100001000100001000100001",  --  5.2939606 -  5.2959084
     "00010000100010000100010000100010",  --  5.2959712 -  5.2979190
     "00010001000100001000100001000100",  --  5.2979819 -  5.2999296
     "00100010000100010000100010000100",  --  5.2999925 -  5.3019403
     "01000010001000010001000100001000",  --  5.3020031 -  5.3039509
     "10000100010000100010000100010000",  --  5.3040137 -  5.3059615
     "10001000100001000100001000100001",  --  5.3060243 -  5.3079721
     "00010000100010001000010001000010",  --  5.3080349 -  5.3099827
     "00100001000100010000100010000100",  --  5.3100456 -  5.3119934
     "01000010001000100001000100001000",  --  5.3120562 -  5.3140040
     "10000100010001000010001000010001",  --  5.3140668 -  5.3160146
     "00010000100010000100010001000010",  --  5.3160774 -  5.3180252
     "00100001000100010000100010000100",  --  5.3180880 -  5.3200358
     "01000100001000100001000100010000",  --  5.3200987 -  5.3220465
     "10001000010001000100001000100001",  --  5.3221093 -  5.3240571
     "00010001000010001000100001000100",  --  5.3241199 -  5.3260677
     "00100010001000010001000100001000",  --  5.3261305 -  5.3280783
     "10000100010001000010001000100001",  --  5.3281411 -  5.3300889
     "00010001000010001000100001000100",  --  5.3301518 -  5.3320995
     "00100010001000010001000100001000",  --  5.3321624 -  5.3341102
     "10001000010001000100001000100010",  --  5.3341730 -  5.3361208
     "00010001000100001000100010000100",  --  5.3361836 -  5.3381314
     "01000100001000100010000100010001",  --  5.3381942 -  5.3401420
     "00001000100010000100010001000010",  --  5.3402049 -  5.3421526
     "00100010000100010001000100001000",  --  5.3422155 -  5.3441633
     "10001000010001000100001000100010",  --  5.3442261 -  5.3461739
     "00010001000100010000100010001000",  --  5.3462367 -  5.3481845
     "01000100010001000010001000100001",  --  5.3482473 -  5.3501951
     "00010001000100001000100010000100",  --  5.3502580 -  5.3522057
     "01000100010000100010001000010001",  --  5.3522686 -  5.3542164
     "00010001000010001000100010000100",  --  5.3542792 -  5.3562270
     "01000100010000100010001000010001",  --  5.3562898 -  5.3582376
     "00010001000010001000100010000100",  --  5.3583004 -  5.3602482
     "01000100010000100010001000100001",  --  5.3603110 -  5.3622588
     "00010001000100001000100010001000",  --  5.3623217 -  5.3642695
     "10000100010001000100001000100010",  --  5.3643323 -  5.3662801
     "00100001000100010001000100001000",  --  5.3663429 -  5.3682907
     "10001000100001000100010001000100",  --  5.3683535 -  5.3703013
     "00100010001000100010000100010001",  --  5.3703641 -  5.3723119
     "00010000100010001000100010000100",  --  5.3723748 -  5.3743226
     "01000100010001000010001000100010",  --  5.3743854 -  5.3763332
     "00100010000100010001000100010000",  --  5.3763960 -  5.3783438
     "10001000100010001000010001000100",  --  5.3784066 -  5.3803544
     "01000100010000100010001000100010",  --  5.3804172 -  5.3823650
     "00100001000100010001000100010000",  --  5.3824279 -  5.3843756
     "10001000100010001000100001000100",  --  5.3844385 -  5.3863863
     "01000100010001000010001000100010",  --  5.3864491 -  5.3883969
     "00100010001000010001000100010001",  --  5.3884597 -  5.3904075
     "00010001000010001000100010001000",  --  5.3904703 -  5.3924181
     "10001000010001000100010001000100",  --  5.3924810 -  5.3944287
     "01000100001000100010001000100010",  --  5.3944916 -  5.3964394
     "00100010000100010001000100010001",  --  5.3965022 -  5.3984500
     "00010001000100001000100010001000",  --  5.3985128 -  5.4004606
     "10001000100010001000100001000100",  --  5.4005234 -  5.4024712
     "01000100010001000100010001000100",  --  5.4025341 -  5.4044818
     "00100010001000100010001000100010",  --  5.4045447 -  5.4064925
     "00100010001000100001000100010001",  --  5.4065553 -  5.4085031
     "00010001000100010001000100010001",  --  5.4085659 -  5.4105137
     "00010000100010001000100010001000",  --  5.4105765 -  5.4125243
     "10001000100010001000100010001000",  --  5.4125872 -  5.4145349
     "10001000010001000100010001000100",  --  5.4145978 -  5.4165456
     "01000100010001000100010001000100",  --  5.4166084 -  5.4185562
     "01000100010001000100010001000100",  --  5.4186190 -  5.4205668
     "00100010001000100010001000100010",  --  5.4206296 -  5.4225774
     "00100010001000100010001000100010",  --  5.4226402 -  5.4245880
     "00100010001000100010001000100010",  --  5.4246509 -  5.4265987
     "00100010001000100010001000100010",  --  5.4266615 -  5.4286093
     "00100010001000100010001000100010",  --  5.4286721 -  5.4306199
     "00100010001000100010001000100010",  --  5.4306827 -  5.4326305
     "00100010001000100010001000100010",  --  5.4326933 -  5.4346411
     "00100010001000100010001000100010",  --  5.4347040 -  5.4366518
     "00100010001000100010001000100010",  --  5.4367146 -  5.4386624
     "00100010001000100010001000100100",  --  5.4387252 -  5.4406730
     "01000100010001000100010001000100",  --  5.4407358 -  5.4426836
     "01000100010001000100010001000100",  --  5.4427464 -  5.4446942
     "01000100010001000100010010001000",  --  5.4447571 -  5.4467048
     "10001000100010001000100010001000",  --  5.4467677 -  5.4487155
     "10001000100010001000100100010001",  --  5.4487783 -  5.4507261
     "00010001000100010001000100010001",  --  5.4507889 -  5.4527367
     "00010001000100100010001000100010",  --  5.4527995 -  5.4547473
     "00100010001000100010001000100100",  --  5.4548102 -  5.4567579
     "01000100010001000100010001000100",  --  5.4568208 -  5.4587686
     "01001000100010001000100010001000",  --  5.4588314 -  5.4607792
     "10001000100100010001000100010001",  --  5.4608420 -  5.4627898
     "00010001000100100010001000100010",  --  5.4628526 -  5.4648004
     "00100010001001000100010001000100",  --  5.4648633 -  5.4668110
     "01000100010010001000100010001000",  --  5.4668739 -  5.4688217
     "10001000100100010001000100010001",  --  5.4688845 -  5.4708323
     "00010010001000100010001000100010",  --  5.4708951 -  5.4728429
     "01000100010001000100010001001000",  --  5.4729057 -  5.4748535
     "10001000100010001000100100010001",  --  5.4749163 -  5.4768641
     "00010001000100100010001000100010",  --  5.4769270 -  5.4788748
     "00100100010001000100010001001000",  --  5.4789376 -  5.4808854
     "10001000100010001001000100010001",  --  5.4809482 -  5.4828960
     "00010010001000100010001000100100",  --  5.4829588 -  5.4849066
     "01000100010001001000100010001000",  --  5.4849694 -  5.4869172
     "10010001000100010001001000100010",  --  5.4869801 -  5.4889279
     "00100010010001000100010001001000",  --  5.4889907 -  5.4909385
     "10001000100010010001000100010001",  --  5.4910013 -  5.4929491
     "00100010001000100100010001000100",  --  5.4930119 -  5.4949597
     "01001000100010001001000100010001",  --  5.4950225 -  5.4969703
     "00010010001000100010010001000100",  --  5.4970332 -  5.4989809
     "01001000100010001000100100010001",  --  5.4990438 -  5.5009916
     "00010010001000100010010001000100",  --  5.5010544 -  5.5030022
     "01001000100010001001000100010001",  --  5.5030650 -  5.5050128
     "00100010001000100100010001000100",  --  5.5050756 -  5.5070234
     "10001000100010010001000100100010",  --  5.5070863 -  5.5090340
     "00100010010001000100010010001000",  --  5.5090969 -  5.5110447
     "10010001000100010010001000100010",  --  5.5111075 -  5.5130553
     "01000100010010001000100010010001",  --  5.5131181 -  5.5150659
     "00010010001000100010010001000100",  --  5.5151287 -  5.5170765
     "10001000100100010001000100100010",  --  5.5171394 -  5.5190871
     "00100100010001001000100010001001",  --  5.5191500 -  5.5210978
     "00010001001000100010010001000100",  --  5.5211606 -  5.5231084
     "10001000100010010001000100100010",  --  5.5231712 -  5.5251190
     "00100100010001001000100010010001",  --  5.5251818 -  5.5271296
     "00010010001000100100010001001000",  --  5.5271925 -  5.5291402
     "10001001000100010010001000100100",  --  5.5292031 -  5.5311509
     "01000100100010001001000100010010",  --  5.5312137 -  5.5331615
     "00100010010001000100100010001001",  --  5.5332243 -  5.5351721
     "00010010001000100100010001001000",  --  5.5352349 -  5.5371827
     "10001001000100010010001001000100",  --  5.5372455 -  5.5391933
     "01001000100010010001001000100010",  --  5.5392562 -  5.5412040
     "01000100010010001001000100010010",  --  5.5412668 -  5.5432146
     "00100010010001001000100010010001",  --  5.5432774 -  5.5452252
     "00010010001001000100010010001001",  --  5.5452880 -  5.5472358
     "00010001001000100100010001001000",  --  5.5472986 -  5.5492464
     "10010001000100100010010001000100",  --  5.5493093 -  5.5512571
     "10001001000100010010001001000100",  --  5.5513199 -  5.5532677
     "01001000100100010001001000100100",  --  5.5533305 -  5.5552783
     "01001000100010010001001000100010",  --  5.5553411 -  5.5572889
     "01000100100010010001000100100010",  --  5.5573517 -  5.5592995
     "01000100100010010001000100100010",  --  5.5593624 -  5.5613101
     "01000100100010001001000100100010",  --  5.5613730 -  5.5633208
     "01000100100010001001000100100010",  --  5.5633836 -  5.5653314
     "01000100100010001001000100100010",  --  5.5653942 -  5.5673420
     "01000100100010010001000100100010",  --  5.5674048 -  5.5693526
     "01000100100010010001001000100100",  --  5.5694155 -  5.5713632
     "01001000100010010001001000100100",  --  5.5714261 -  5.5733739
     "01001000100100010010001001000100",  --  5.5734367 -  5.5753845
     "10001001000100100010001001000100",  --  5.5754473 -  5.5773951
     "10001001000100100010010001001000",  --  5.5774579 -  5.5794057
     "10010001001000100100010010001001",  --  5.5794686 -  5.5814163
     "00010010001001000100100010010001",  --  5.5814792 -  5.5834270
     "00100010010001001000100100010010",  --  5.5834898 -  5.5854376
     "00100100010010001001001000100100",  --  5.5855004 -  5.5874482
     "01001000100100010010001001000100",  --  5.5875110 -  5.5894588
     "10001001000100100010010001001001",  --  5.5895216 -  5.5914694
     "00010010001001000100100010010001",  --  5.5915323 -  5.5934801
     "00100010010001001001000100100010",  --  5.5935429 -  5.5954907
     "01000100100010010001001001000100",  --  5.5955535 -  5.5975013
     "10001001000100100010010001001001",  --  5.5975641 -  5.5995119
     "00010010001001000100100100010010",  --  5.5995747 -  5.6015225
     "00100100010010001001001000100100",  --  5.6015854 -  5.6035332
     "01001000100100100010010001001000",  --  5.6035960 -  5.6055438
     "10010010001001000100100010010010",  --  5.6056066 -  5.6075544
     "00100100010010010001001000100100",  --  5.6076172 -  5.6095650
     "01001001000100100010010010001001",  --  5.6096278 -  5.6115756
     "00010010001001001000100100010010",  --  5.6116385 -  5.6135862
     "01000100100010010010001001000100",  --  5.6136491 -  5.6155969
     "10010001001001000100100010010010",  --  5.6156597 -  5.6176075
     "00100100010010010001001000100100",  --  5.6176703 -  5.6196181
     "10001001001000100100010010010001",  --  5.6196809 -  5.6216287
     "00100010010010001001001000100100",  --  5.6216916 -  5.6236393
     "01001001000100100100010010010001",  --  5.6237022 -  5.6256500
     "00100010010010001001001000100100",  --  5.6257128 -  5.6276606
     "10001001000100100100010010010001",  --  5.6277234 -  5.6296712
     "00100100010010010001001001000100",  --  5.6297340 -  5.6316818
     "10001001001000100100100010010010",  --  5.6317447 -  5.6336924
     "00100100100010010010001001001000",  --  5.6337553 -  5.6357031
     "10010010001001001000100100100010",  --  5.6357659 -  5.6377137
     "01001000100100100010010010001001",  --  5.6377765 -  5.6397243
     "00100010010010001001001000100100",  --  5.6397871 -  5.6417349
     "10010001001001000100100100010010",  --  5.6417978 -  5.6437455
     "01000100100100010010010010001001",  --  5.6438084 -  5.6457562
     "00100010010010001001001000100100",  --  5.6458190 -  5.6477668
     "10010001001001000100100100010010",  --  5.6478296 -  5.6497774
     "01001000100100100010010010010001",  --  5.6498402 -  5.6517880
     "00100100010010010010001001001000",  --  5.6518508 -  5.6537986
     "10010010010001001001000100100100",  --  5.6538615 -  5.6558093
     "10001001001000100100100100010010",  --  5.6558721 -  5.6578199
     "01001000100100100010010010010001",  --  5.6578827 -  5.6598305
     "00100100100010010010010001001001",  --  5.6598933 -  5.6618411
     "00100010010010010001001001000100",  --  5.6619039 -  5.6638517
     "10010010001001001001000100100100",  --  5.6639146 -  5.6658624
     "10001001001001000100100100100010",  --  5.6659252 -  5.6678730
     "01001001001000100100100100010010",  --  5.6679358 -  5.6698836
     "01001000100100100100010010010010",  --  5.6699464 -  5.6718942
     "01000100100100100010010010010001",  --  5.6719570 -  5.6739048
     "00100100100100010010010010001001",  --  5.6739677 -  5.6759154
     "00100100100010010010010001001001",  --  5.6759783 -  5.6779261
     "00100100010010010010010001001001",  --  5.6779889 -  5.6799367
     "00100100010010010010001001001001",  --  5.6799995 -  5.6819473
     "00100010010010010010001001001001",  --  5.6820101 -  5.6839579
     "00100010010010010010010001001001",  --  5.6840208 -  5.6859685
     "00100100010010010010010001001001",  --  5.6860314 -  5.6879792
     "00100100010010010010010010001001",  --  5.6880420 -  5.6899898
     "00100100100010010010010010010001",  --  5.6900526 -  5.6920004
     "00100100100100100010010010010010",  --  5.6920632 -  5.6940110
     "01000100100100100100100010010010",  --  5.6940739 -  5.6960216
     "01001001000100100100100100100010",  --  5.6960845 -  5.6980323
     "01001001001001000100100100100100",  --  5.6980951 -  5.7000429
     "10010001001001001001001000100100",  --  5.7001057 -  5.7020535
     "10010010010010001001001001001001",  --  5.7021163 -  5.7040641
     "00100010010010010010010010010001",  --  5.7041269 -  5.7060747
     "00100100100100100100010010010010",  --  5.7061376 -  5.7080854
     "01001001001000100100100100100100",  --  5.7081482 -  5.7100960
     "10001001001001001001001001001000",  --  5.7101588 -  5.7121066
     "10010010010010010010010001001001",  --  5.7121694 -  5.7141172
     "00100100100100100100010010010010",  --  5.7141800 -  5.7161278
     "01001001001001000100100100100100",  --  5.7161907 -  5.7181385
     "10010010010010001001001001001001",  --  5.7182013 -  5.7201491
     "00100100100100010010010010010010",  --  5.7202119 -  5.7221597
     "01001001001001000100100100100100",  --  5.7222225 -  5.7241703
     "10010010010010010001001001001001",  --  5.7242331 -  5.7261809
     "00100100100100100100100100010010",  --  5.7262438 -  5.7281915
     "01001001001001001001001001001001",  --  5.7282544 -  5.7302022
     "00010010010010010010010010010010",  --  5.7302650 -  5.7322128
     "01001001001001000100100100100100",  --  5.7322756 -  5.7342234
     "10010010010010010010010010010010",  --  5.7342862 -  5.7362340
     "01000100100100100100100100100100",  --  5.7362969 -  5.7382446
     "10010010010010010010010010010010",  --  5.7383075 -  5.7402553
     "00100100100100100100100100100100",  --  5.7403181 -  5.7422659
     "10010010010010010010010010010010",  --  5.7423287 -  5.7442765
     "01001001001001001000100100100100",  --  5.7443393 -  5.7462871
     "10010010010010010010010010010010",  --  5.7463500 -  5.7482977
     "01001001001001001001001001001001",  --  5.7483606 -  5.7503084
     "00100100100100100100100100100100",  --  5.7503712 -  5.7523190
     "10010010010010010010010010010010",  --  5.7523818 -  5.7543296
     "01001001001001001001001001001001",  --  5.7543924 -  5.7563402
     "00100100100100100100100100100100",  --  5.7564031 -  5.7583508
     "10010010010010010010010010010010",  --  5.7584137 -  5.7603615
     "01001001001001001001001001001001",  --  5.7604243 -  5.7623721
     "00100100100100100100100100100100",  --  5.7624349 -  5.7643827
     "10010010010010010010010010010010",  --  5.7644455 -  5.7663933
     "01001001001001001001001001001001",  --  5.7664561 -  5.7684039
     "00100100101001001001001001001001",  --  5.7684668 -  5.7704146
     "00100100100100100100100100100100",  --  5.7704774 -  5.7724252
     "10010010010010010010010010100100",  --  5.7724880 -  5.7744358
     "10010010010010010010010010010010",  --  5.7744986 -  5.7764464
     "01001001001001001001001010010010",  --  5.7765092 -  5.7784570
     "01001001001001001001001001001001",  --  5.7785199 -  5.7804677
     "00100100100101001001001001001001",  --  5.7805305 -  5.7824783
     "00100100100100100100100101001001",  --  5.7825411 -  5.7844889
     "00100100100100100100100100100100",  --  5.7845517 -  5.7864995
     "10100100100100100100100100100100",  --  5.7865623 -  5.7885101
     "10010010100100100100100100100100",  --  5.7885730 -  5.7905207
     "10010010010100100100100100100100",  --  5.7905836 -  5.7925314
     "10010010010100100100100100100100",  --  5.7925942 -  5.7945420
     "10010010010100100100100100100100",  --  5.7946048 -  5.7965526
     "10010010100100100100100100100100",  --  5.7966154 -  5.7985632
     "10010100100100100100100100100101",  --  5.7986261 -  5.8005738
     "00100100100100100100100101001001",  --  5.8006367 -  5.8025845
     "00100100100100100101001001001001",  --  5.8026473 -  5.8045951
     "00100100101001001001001001001001",  --  5.8046579 -  5.8066057
     "00101001001001001001001001010010",  --  5.8066685 -  5.8086163
     "01001001001001010010010010010010",  --  5.8086792 -  5.8106269
     "01001010010010010010010010100100",  --  5.8106898 -  5.8126376
     "10010010010010100100100100100100",  --  5.8127004 -  5.8146482
     "10100100100100100100101001001001",  --  5.8147110 -  5.8166588
     "00100100101001001001001001001010",  --  5.8167216 -  5.8186694
     "01001001001001010010010010010010",  --  5.8187322 -  5.8206800
     "01010010010010010010100100100100",  --  5.8207429 -  5.8226907
     "10010100100100100100101001001001",  --  5.8227535 -  5.8247013
     "00100101001001001001001010010010",  --  5.8247641 -  5.8267119
     "01001001010010010010010100100100",  --  5.8267747 -  5.8287225
     "10010010100100100100100101001001",  --  5.8287853 -  5.8307331
     "00100101001001001001001010010010",  --  5.8307960 -  5.8327438
     "01001010010010010010100100100100",  --  5.8328066 -  5.8347544
     "10100100100100100101001001001001",  --  5.8348172 -  5.8367650
     "01001001001001010010010010010100",  --  5.8368278 -  5.8387756
     "10010010010100100100100101001001",  --  5.8388384 -  5.8407862
     "00100101001001001010010010010010",  --  5.8408491 -  5.8427968
     "10010010010010100100100100101001",  --  5.8428597 -  5.8448075
     "00100101001001001001010010010010",  --  5.8448703 -  5.8468181
     "10010010010010100100100101001001",  --  5.8468809 -  5.8488287
     "00100101001001001010010010010010",  --  5.8488915 -  5.8508393
     "10010010010100100100101001001001",  --  5.8509022 -  5.8528499
     "00101001001001010010010010100100",  --  5.8529128 -  5.8548606
     "10010100100100100101001001001010",  --  5.8549234 -  5.8568712
     "01001001010010010010100100100101",  --  5.8569340 -  5.8588818
     "00100100101001001001010010010010",  --  5.8589446 -  5.8608924
     "10010010010100100100101001001001",  --  5.8609553 -  5.8629030
     "01001001001010010010100100100101",  --  5.8629659 -  5.8649137
     "00100100101001001001010010010010",  --  5.8649765 -  5.8669243
     "10010010100100100101001001001010",  --  5.8669871 -  5.8689349
     "01001001010010010100100100101001",  --  5.8689977 -  5.8709455
     "00100101001001010010010010100100",  --  5.8710084 -  5.8729561
     "10100100100101001001010010010010",  --  5.8730190 -  5.8749668
     "10010010100100100101001001010010",  --  5.8750296 -  5.8769774
     "01001010010010100100100101001001",  --  5.8770402 -  5.8789880
     "01001001001010010010100100101001",  --  5.8790508 -  5.8809986
     "00100101001001010010010100100100",  --  5.8810614 -  5.8830092
     "10100100101001001010010010010100",  --  5.8830721 -  5.8850199
     "10010100100101001001010010010010",  --  5.8850827 -  5.8870305
     "10010010100100101001001010010010",  --  5.8870933 -  5.8890411
     "10010010100100100101001001010010",  --  5.8891039 -  5.8910517
     "01010010010100100101001001010010",  --  5.8911145 -  5.8930623
     "01010010010100100101001001001010",  --  5.8931252 -  5.8950730
     "01001010010010100100101001001010",  --  5.8951358 -  5.8970836
     "01001010010010100100101001001010",  --  5.8971464 -  5.8990942
     "01001010010100100101001001010010",  --  5.8991570 -  5.9011048
     "01010010010100100101001001010010",  --  5.9011676 -  5.9031154
     "01010010010100100101001001010010",  --  5.9031783 -  5.9051260
     "10010010100100101001001010010010",  --  5.9051889 -  5.9071367
     "10010010100101001001010010010100",  --  5.9071995 -  5.9091473
     "10010100101001001010010010100100",  --  5.9092101 -  5.9111579
     "10100101001001010010010100100101",  --  5.9112207 -  5.9131685
     "00101001001010010010100100101001",  --  5.9132314 -  5.9151791
     "01001001010010010100101001001010",  --  5.9152420 -  5.9171898
     "01001010010100100101001010010010",  --  5.9172526 -  5.9192004
     "10010010100101001001010010010100",  --  5.9192632 -  5.9212110
     "10100100101001010010010100101001",  --  5.9212738 -  5.9232216
     "00101001001010010100100101001010",  --  5.9232845 -  5.9252322
     "01001010010100100101001010010010",  --  5.9252951 -  5.9272429
     "10010100100101001010010010100101",  --  5.9273057 -  5.9292535
     "00100101001010010010100101001001",  --  5.9293163 -  5.9312641
     "01001010010010100101001001010010",  --  5.9313269 -  5.9332747
     "10010100100101001010010010100101",  --  5.9333375 -  5.9352853
     "00100101001010010100100101001010",  --  5.9353482 -  5.9372960
     "01001010010100101001001010010100",  --  5.9373588 -  5.9393066
     "10100100101001010010100100101001",  --  5.9393694 -  5.9413172
     "01001010010010100101001010010010",  --  5.9413800 -  5.9433278
     "10010100101001001010010100101001",  --  5.9433906 -  5.9453384
     "00101001010010100101001001010010",  --  5.9454013 -  5.9473491
     "10010100100101001010010100101001",  --  5.9474119 -  5.9493597
     "00101001010010100101001001010010",  --  5.9494225 -  5.9513703
     "10010100101001010010010100101001",  --  5.9514331 -  5.9533809
     "01001010010010100101001010010100",  --  5.9534437 -  5.9553915
     "10100100101001010010100101001010",  --  5.9554544 -  5.9574021
     "01010010010100101001010010100101",  --  5.9574650 -  5.9594128
     "00101001001010010100101001010010",  --  5.9594756 -  5.9614234
     "10010100101001010010010100101001",  --  5.9614862 -  5.9634340
     "01001010010100101001010010100100",  --  5.9634968 -  5.9654446
     "10100101001010010100101001010010",  --  5.9655075 -  5.9674552
     "10010100101001010010100101001010",  --  5.9675181 -  5.9694659
     "01001010010100101001010010100101",  --  5.9695287 -  5.9714765
     "00101001010010100101001010010100",  --  5.9715393 -  5.9734871
     "10100101001010010100101001010010",  --  5.9735499 -  5.9754977
     "10010100101001010010100101001010",  --  5.9755606 -  5.9775083
     "01010010100101001010010100101001",  --  5.9775712 -  5.9795190
     "01001010010100101001010010100101",  --  5.9795818 -  5.9815296
     "00101001010010100101001010010100",  --  5.9815924 -  5.9835402
     "10100101001010010100101010010100",  --  5.9836030 -  5.9855508
     "10100101001010010100101001010010",  --  5.9856137 -  5.9875614
     "10010100101001010010100101010010",  --  5.9876243 -  5.9895721
     "10010100101001010010100101001010",  --  5.9896349 -  5.9915827
     "01010010101001010010100101001010",  --  5.9916455 -  5.9935933
     "01010010100101010010100101001010",  --  5.9936561 -  5.9956039
     "01010010100101001010100101001010",  --  5.9956667 -  5.9976145
     "01010010100101010010100101001010",  --  5.9976774 -  5.9996252
     "01010010100101010010100101001010",  --  5.9996880 -  6.0016358
     "01010010101001010010100101001010",  --  6.0016986 -  6.0036464
     "10010100101001010010101001010010",  --  6.0037092 -  6.0056570
     "10010100101010010100101001010010",  --  6.0057198 -  6.0076676
     "10100101001010010100101010010100",  --  6.0077305 -  6.0096783
     "10100101010010100101001010010101",  --  6.0097411 -  6.0116889
     "00101001010010101001010010100101",  --  6.0117517 -  6.0136995
     "01001010010100101010010100101001",  --  6.0137623 -  6.0157101
     "01010010100101001010100101001010",  --  6.0157729 -  6.0177207
     "10010100101001010100101001010010",  --  6.0177836 -  6.0197313
     "10100101001010100101001010010101",  --  6.0197942 -  6.0217420
     "00101001010100101001010100101001",  --  6.0218048 -  6.0237526
     "01001010100101001010100101001010",  --  6.0238154 -  6.0257632
     "10010100101010010100101010010100",  --  6.0258260 -  6.0277738
     "10100101010010100101010010100101",  --  6.0278367 -  6.0297844
     "01001010010101001010100101001010",  --  6.0298473 -  6.0317951
     "10010100101010010100101010010100",  --  6.0318579 -  6.0338057
     "10101001010010101001010010101001",  --  6.0338685 -  6.0358163
     "01010010100101010010100101010010",  --  6.0358791 -  6.0378269
     "10100101001010100101001010100101",  --  6.0378898 -  6.0398375
     "01001010010101001010100101001010",  --  6.0399004 -  6.0418482
     "10010101001010010101001010100101",  --  6.0419110 -  6.0438588
     "00101010010101001010010101001010",  --  6.0439216 -  6.0458694
     "10010100101010010101001010010101",  --  6.0459322 -  6.0478800
     "00101010010101001010010101001010",  --  6.0479428 -  6.0498906
     "10010101001010010101001010100101",  --  6.0499535 -  6.0519013
     "01001010100101001010100101010010",  --  6.0519641 -  6.0539119
     "10100101010010100101010010101001",  --  6.0539747 -  6.0559225
     "01010010101001010100101010010100",  --  6.0559853 -  6.0579331
     "10101001010100101010010101001010",  --  6.0579959 -  6.0599437
     "10010101001010100101010010101001",  --  6.0600066 -  6.0619544
     "01001010100101010010101001010100",  --  6.0620172 -  6.0639650
     "10101001010100101010010101001010",  --  6.0640278 -  6.0659756
     "10010101001010100101010010101001",  --  6.0660384 -  6.0679862
     "01010010101001010100101010010101",  --  6.0680490 -  6.0699968
     "00101010010101010010101001010100",  --  6.0700597 -  6.0720074
     "10101001010100101010010101001010",  --  6.0720703 -  6.0740181
     "10010101001010101001010100101010",  --  6.0740809 -  6.0760287
     "01010100101010010101001010101001",  --  6.0760915 -  6.0780393
     "01010010101001010100101010010101",  --  6.0781021 -  6.0800499
     "01001010100101010010101001010101",  --  6.0801128 -  6.0820605
     "00101010010101001010100101010100",  --  6.0821234 -  6.0840712
     "10101001010100101010100101010010",  --  6.0841340 -  6.0860818
     "10100101010100101010010101001010",  --  6.0861446 -  6.0880924
     "10100101010010101010010101001010",  --  6.0881552 -  6.0901030
     "10010101010010101001010101001010",  --  6.0901659 -  6.0921136
     "10010101010010101001010101001010",  --  6.0921765 -  6.0941243
     "10010101010010101001010101001010",  --  6.0941871 -  6.0961349
     "10010101010010101010010101001010",  --  6.0961977 -  6.0981455
     "10100101010010101010010101010010",  --  6.0982083 -  6.1001561
     "10100101010100101010010101010010",  --  6.1002190 -  6.1021667
     "10101001010101001010100101010100",  --  6.1022296 -  6.1041774
     "10101010010101001010101001010101",  --  6.1042402 -  6.1061880
     "00101010100101010100101010010101",  --  6.1062508 -  6.1081986
     "01001010101001010101001010101001",  --  6.1082614 -  6.1102092
     "01010100101010100101010010101010",  --  6.1102720 -  6.1122198
     "01010101001010101001010101001010",  --  6.1122827 -  6.1142305
     "10100101010100101010100101010100",  --  6.1142933 -  6.1162411
     "10101010010101010010101010010101",  --  6.1163039 -  6.1182517
     "01001010101010010101010010101010",  --  6.1183145 -  6.1202623
     "01010101001010101001010101001010",  --  6.1203251 -  6.1222729
     "10100101010101001010101001010101",  --  6.1223358 -  6.1242836
     "00101010100101010101001010101001",  --  6.1243464 -  6.1262942
     "01010100101010101001010101001010",  --  6.1263570 -  6.1283048
     "10100101010101001010101001010101",  --  6.1283676 -  6.1303154
     "01001010101001010101010010101010",  --  6.1303782 -  6.1323260
     "01010101010010101010010101010100",  --  6.1323889 -  6.1343366
     "10101010010101010100101010101001",  --  6.1343995 -  6.1363473
     "01010100101010101001010101010010",  --  6.1364101 -  6.1383579
     "10101001010101010010101010100101",  --  6.1384207 -  6.1403685
     "01010100101010101001010101001010",  --  6.1404313 -  6.1423791
     "10101001010101010010101010100101",  --  6.1424420 -  6.1443897
     "01010100101010101001010101010010",  --  6.1444526 -  6.1464004
     "10101010010101010100101010101001",  --  6.1464632 -  6.1484110
     "01010101001010101010010101010100",  --  6.1484738 -  6.1504216
     "10101010101001010101010010101010",  --  6.1504844 -  6.1524322
     "10010101010101001010101010010101",  --  6.1524951 -  6.1544428
     "01010010101010101001010101010010",  --  6.1545057 -  6.1564535
     "10101010100101010101001010101010",  --  6.1565163 -  6.1584641
     "10010101010100101010101010010101",  --  6.1585269 -  6.1604747
     "01010010101010101001010101010100",  --  6.1605375 -  6.1624853
     "10101010101001010101010010101010",  --  6.1625481 -  6.1644959
     "10100101010101010010101010101001",  --  6.1645588 -  6.1665066
     "01010101010010101010101001010101",  --  6.1665694 -  6.1685172
     "01010010101010101001010101010100",  --  6.1685800 -  6.1705278
     "10101010101010010101010101001010",  --  6.1705906 -  6.1725384
     "10101010010101010101010010101010",  --  6.1726012 -  6.1745490
     "10100101010101010100101010101010",  --  6.1746119 -  6.1765597
     "01010101010101001010101010100101",  --  6.1766225 -  6.1785703
     "01010101010010101010101010010101",  --  6.1786331 -  6.1805809
     "01010101001010101010101001010101",  --  6.1806437 -  6.1825915
     "01010100101010101010100101010101",  --  6.1826543 -  6.1846021
     "01010010101010101010010101010101",  --  6.1846650 -  6.1866127
     "01001010101010101010010101010101",  --  6.1866756 -  6.1886234
     "01001010101010101010010101010101",  --  6.1886862 -  6.1906340
     "01001010101010101010010101010101",  --  6.1906968 -  6.1926446
     "01010010101010101010100101010101",  --  6.1927074 -  6.1946552
     "01010100101010101010101001010101",  --  6.1947181 -  6.1966658
     "01010101001010101010101010100101",  --  6.1967287 -  6.1986765
     "01010101010100101010101010101001",  --  6.1987393 -  6.2006871
     "01010101010101010010101010101010",  --  6.2007499 -  6.2026977
     "10100101010101010101010010101010",  --  6.2027605 -  6.2047083
     "10101010100101010101010101010010",  --  6.2047712 -  6.2067189
     "10101010101010101001010101010101",  --  6.2067818 -  6.2087296
     "01010010101010101010101010010101",  --  6.2087924 -  6.2107402
     "01010101010101001010101010101010",  --  6.2108030 -  6.2127508
     "10100101010101010101010101001010",  --  6.2128136 -  6.2147614
     "10101010101010100101010101010101",  --  6.2148243 -  6.2167720
     "01010100101010101010101010101001",  --  6.2168349 -  6.2187827
     "01010101010101010101001010101010",  --  6.2188455 -  6.2207933
     "10101010101010010101010101010101",  --  6.2208561 -  6.2228039
     "01010100101010101010101010101010",  --  6.2228667 -  6.2248145
     "01010101010101010101010101001010",  --  6.2248773 -  6.2268251
     "10101010101010101010100101010101",  --  6.2268880 -  6.2288358
     "01010101010101010010101010101010",  --  6.2288986 -  6.2308464
     "10101010101010010101010101010101",  --  6.2309092 -  6.2328570
     "01010101010010101010101010101010",  --  6.2329198 -  6.2348676
     "10101010100101010101010101010101",  --  6.2349304 -  6.2368782
     "01010101010010101010101010101010",  --  6.2369411 -  6.2388889
     "10101010101001010101010101010101",  --  6.2389517 -  6.2408995
     "01010101010101010010101010101010",  --  6.2409623 -  6.2429101
     "10101010101010101010100101010101",  --  6.2429729 -  6.2449207
     "01010101010101010101010101010010",  --  6.2449835 -  6.2469313
     "10101010101010101010101010101010",  --  6.2469942 -  6.2489419
     "10101010100101010101010101010101",  --  6.2490048 -  6.2509526
     "01010101010101010101010010101010",  --  6.2510154 -  6.2529632
     "10101010101010101010101010101010",  --  6.2530260 -  6.2549738
     "10101010101001010101010101010101",  --  6.2550366 -  6.2569844
     "01010101010101010101010101010101",  --  6.2570473 -  6.2589950
     "01010100101010101010101010101010",  --  6.2590579 -  6.2610057
     "10101010101010101010101010101010",  --  6.2610685 -  6.2630163
     "10101010101001010101010101010101",  --  6.2630791 -  6.2650269
     "01010101010101010101010101010101",  --  6.2650897 -  6.2670375
     "01010101010101010101010101010101",  --  6.2671004 -  6.2690481
     "01010100101010101010101010101010",  --  6.2691110 -  6.2710588
     "10101010101010101010101010101010",  --  6.2711216 -  6.2730694
     "10101010101010101010101010101010",  --  6.2731322 -  6.2750800
     "10101010101010101010101010101010",  --  6.2751428 -  6.2770906
     "10101010101010101010101010101010",  --  6.2771534 -  6.2791012
     "10101010101010101010101010101010",  --  6.2791641 -  6.2811119
     "10101010101010101010101010101010"); --  6.2811747 -  6.2831225
begin

process(clk100MHz)
    begin
        if rising_edge(clK100MHz) then
            if (mask and data) = x"00000000" then
                pin <= '0';
            else
                pin <= '1';
            end if;

            data <= memory(to_integer(addr));

            mask <= mask(30 downto 0) & mask(31); 
            if mask(30) = '1' then
                if addr = memory'high then
                    addr <= (others => '0');
                else
                    addr <= addr + 1;
                end if;
            end if;
        end if;
    end process;
end whatever;
